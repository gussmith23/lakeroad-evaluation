module uge2_2(input  [1:0] a, input  [1:0] b, output  out);
  assign out = a >= b;
endmodule
