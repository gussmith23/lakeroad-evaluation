module uge7_2(input unsigned[6:0] a, input unsigned[6:0] b, output unsigned out);
  assign out = a >= b;
endmodule
