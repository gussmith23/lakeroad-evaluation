module example(input [15:0] a, output [0:0] out);
  assign out = a[15];
endmodule
