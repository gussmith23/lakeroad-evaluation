module sgt3_2(input signed [2:0] a, input signed [2:0] b, output signed out);
  assign out = a > b;
endmodule
