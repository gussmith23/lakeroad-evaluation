module not4_1(input  [3:0] a, output [3:0] out);
  assign out = ~a;
endmodule
