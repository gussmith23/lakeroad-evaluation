module ult5_2(input  [4:0] a, input  [4:0] b, output  out);
  assign out = a < b;
endmodule
