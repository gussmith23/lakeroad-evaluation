module parity96_1(input  [95:0] a, output out);
  assign out = ^a;
endmodule
