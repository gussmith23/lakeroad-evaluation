module slt2_2(input signed[1:0] a, input signed[1:0] b, output signed out);
  assign out = a < b;
endmodule
