module ule3_2(input  [2:0] a, input  [2:0] b, output  out);
  assign out = a <= b;
endmodule
