module example(input [7:0] a, output [3:0] out);
  assign out = a[3:0];
endmodule