module ssub5_2(input signed [4:0] a, input signed [4:0] b, output signed[4:0] out);
  assign out = a - b;
endmodule
