module uge7_2(input unsigned[6:0] a, input unsigned[6:0] b, output unsigned[6:0] out);
  assign out = a >= b;
endmodule
