module sadd32_2(input signed [31:0] a, input signed [31:0] b, output signed[31:0] out);
  assign out = a + b;
endmodule
