module divs8_2(input signed[7:0] a, input signed[7:0] b, output signed[7:0] out);
  assign out = a / b;
endmodule
