module ssub64_2(input signed [63:0] a, input signed [63:0] b, output signed[63:0] out);
  assign out = a - b;
endmodule
