module eq8_2(input  [7:0] a, input  [7:0] b, output  out);
  assign out = a == b;
endmodule
