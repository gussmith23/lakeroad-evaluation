module shl3_2(input [2:0] a, input [2:0] b, output [2:0] out);
  assign out = a << b;
endmodule
