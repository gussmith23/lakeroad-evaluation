module extract4_3_0(input [3:0] a, output [2:0] out);
  assign out = a[2:0];
endmodule