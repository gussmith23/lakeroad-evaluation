module ule8_2(input unsigned[7:0] a, input unsigned[7:0] b, output unsigned out);
  assign out = a <= b;
endmodule
