module example(input [7:0] a, output [0:0] out);
  assign out = a[7];
endmodule
