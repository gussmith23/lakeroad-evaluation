/**
 * Core primitives for Calyx.
 * Implements core primitives used by the compiler.
 *
 * Conventions:
 * - All parameter names must be SNAKE_CASE and all caps.
 * - Port names must be snake_case, no caps.
 */
`default_nettype none

module std_const #(
    parameter WIDTH = 32,
    parameter VALUE = 0
) (
   output logic [WIDTH - 1:0] out
);
  assign out = VALUE;
endmodule

module std_wire #(
  parameter WIDTH = 32
) (
  input wire logic [WIDTH - 1:0] in,
  output logic [WIDTH - 1:0] out
);
  assign out = in;
endmodule

module std_slice #(
    parameter IN_WIDTH  = 32,
    parameter OUT_WIDTH = 32
) (
   input wire                   logic [ IN_WIDTH-1:0] in,
   output logic [OUT_WIDTH-1:0] out
);
  assign out = in[OUT_WIDTH-1:0];

  `ifdef VERILATOR
    always_comb begin
      if (IN_WIDTH < OUT_WIDTH)
        $error(
          "std_slice: Input width less than output width\n",
          "IN_WIDTH: %0d", IN_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_pad #(
    parameter IN_WIDTH  = 32,
    parameter OUT_WIDTH = 32
) (
   input wire logic [IN_WIDTH-1:0]  in,
   output logic     [OUT_WIDTH-1:0] out
);
  localparam EXTEND = OUT_WIDTH - IN_WIDTH;
  assign out = { {EXTEND {1'b0}}, in};

  `ifdef VERILATOR
    always_comb begin
      if (IN_WIDTH > OUT_WIDTH)
        $error(
          "std_pad: Output width less than input width\n",
          "IN_WIDTH: %0d", IN_WIDTH,
          "OUT_WIDTH: %0d", OUT_WIDTH
        );
    end
  `endif
endmodule

module std_not #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] in,
   output logic [WIDTH-1:0] out
);
  assign out = ~in;
endmodule

module std_and #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left & right;
endmodule

module std_or #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left | right;
endmodule

module std_xor #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left ^ right;
endmodule

module std_add #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left + right;
endmodule

module std_sub #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module std_gt #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left > right;
endmodule

module std_lt #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left < right;
endmodule

module std_eq #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left == right;
endmodule

module std_neq #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left != right;
endmodule

module std_ge #(
    parameter WIDTH = 32
) (
    input wire   logic [WIDTH-1:0] left,
    input wire   logic [WIDTH-1:0] right,
    output logic out
);
  assign out = left >= right;
endmodule

module std_le #(
    parameter WIDTH = 32
) (
   input wire   logic [WIDTH-1:0] left,
   input wire   logic [WIDTH-1:0] right,
   output logic out
);
  assign out = left <= right;
endmodule

module std_lsh #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left << right;
endmodule

module std_rsh #(
    parameter WIDTH = 32
) (
   input wire               logic [WIDTH-1:0] left,
   input wire               logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
  assign out = left >> right;
endmodule

/// this primitive is intended to be used
/// for lowering purposes (not in source programs)
module std_mux #(
    parameter WIDTH = 32
) (
   input wire               logic cond,
   input wire               logic [WIDTH-1:0] tru,
   input wire               logic [WIDTH-1:0] fal,
   output logic [WIDTH-1:0] out
);
  assign out = cond ? tru : fal;
endmodule

/// Memories
module std_reg #(
    parameter WIDTH = 32
) (
   input wire [ WIDTH-1:0]    in,
   input wire                 write_en,
   input wire                 clk,
   input wire                 reset,
    // output
   output logic [WIDTH - 1:0] out,
   output logic               done
);

  always_ff @(posedge clk) begin
    if (reset) begin
       out <= 0;
       done <= 0;
    end else if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module std_mem_d1 #(
    parameter WIDTH = 32,
    parameter SIZE = 16,
    parameter IDX_SIZE = 4
) (
   input wire                logic [IDX_SIZE-1:0] addr0,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  logic [WIDTH-1:0] mem[SIZE-1:0];

  /* verilator lint_off WIDTH */
  assign read_data = mem[addr0];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0] <= write_data;
      done <= 1'd1;
    end else done <= 1'd0;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= SIZE)
        $error(
          "std_mem_d1: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "SIZE: %0d", SIZE
        );
    end
  `endif
endmodule

module std_mem_d2 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0];

  assign read_data = mem[addr0][addr1];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0][addr1] <= write_data;
      done <= 1'd1;
    end else done <= 1'd0;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d2: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d2: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
    end
  `endif
endmodule

module std_mem_d3 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D2_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4,
    parameter D2_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [D2_IDX_SIZE-1:0] addr2,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0][D2_SIZE-1:0];

  assign read_data = mem[addr0][addr1][addr2];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0][addr1][addr2] <= write_data;
      done <= 1'd1;
    end else done <= 1'd0;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
      if (addr2 >= D2_SIZE)
        $error(
          "std_mem_d3: Out of bounds access\n",
          "addr2: %0d\n", addr2,
          "D2_SIZE: %0d", D2_SIZE
        );
    end
  `endif
endmodule

module std_mem_d4 #(
    parameter WIDTH = 32,
    parameter D0_SIZE = 16,
    parameter D1_SIZE = 16,
    parameter D2_SIZE = 16,
    parameter D3_SIZE = 16,
    parameter D0_IDX_SIZE = 4,
    parameter D1_IDX_SIZE = 4,
    parameter D2_IDX_SIZE = 4,
    parameter D3_IDX_SIZE = 4
) (
   input wire                logic [D0_IDX_SIZE-1:0] addr0,
   input wire                logic [D1_IDX_SIZE-1:0] addr1,
   input wire                logic [D2_IDX_SIZE-1:0] addr2,
   input wire                logic [D3_IDX_SIZE-1:0] addr3,
   input wire                logic [ WIDTH-1:0] write_data,
   input wire                logic write_en,
   input wire                logic clk,
   output logic [ WIDTH-1:0] read_data,
   output logic              done
);

  /* verilator lint_off WIDTH */
  logic [WIDTH-1:0] mem[D0_SIZE-1:0][D1_SIZE-1:0][D2_SIZE-1:0][D3_SIZE-1:0];

  assign read_data = mem[addr0][addr1][addr2][addr3];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0][addr1][addr2][addr3] <= write_data;
      done <= 1'd1;
    end else done <= 1'd0;
  end

  // Check for out of bounds access
  `ifdef VERILATOR
    always_comb begin
      if (addr0 >= D0_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr0: %0d\n", addr0,
          "D0_SIZE: %0d", D0_SIZE
        );
      if (addr1 >= D1_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr1: %0d\n", addr1,
          "D1_SIZE: %0d", D1_SIZE
        );
      if (addr2 >= D2_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr2: %0d\n", addr2,
          "D2_SIZE: %0d", D2_SIZE
        );
      if (addr3 >= D3_SIZE)
        $error(
          "std_mem_d4: Out of bounds access\n",
          "addr3: %0d\n", addr3,
          "D3_SIZE: %0d", D3_SIZE
        );
    end
  `endif
endmodule

`default_nettype wire
module main (
    input logic go,
    input logic clk,
    input logic reset,
    output logic done,
    output logic index_addr0,
    output logic [4:0] index_write_data,
    output logic index_write_en,
    output logic index_clk,
    input logic [4:0] index_read_data,
    input logic index_done
);
    logic tcam_write_en;
    logic tcam_search_en;
    logic [31:0] tcam_in;
    logic [5:0] tcam_prefix_len;
    logic [4:0] tcam_write_index;
    logic [4:0] tcam_index;
    logic tcam_go;
    logic tcam_clk;
    logic tcam_reset;
    logic tcam_done;
    logic [1:0] fsm_in;
    logic fsm_write_en;
    logic fsm_clk;
    logic fsm_reset;
    logic [1:0] fsm_out;
    logic fsm_done;
    logic save_index_go_in;
    logic save_index_go_out;
    logic save_index_done_in;
    logic save_index_done_out;
    logic invoke_go_in;
    logic invoke_go_out;
    logic invoke_done_in;
    logic invoke_done_out;
    logic invoke0_go_in;
    logic invoke0_go_out;
    logic invoke0_done_in;
    logic invoke0_done_out;
    logic tdcc_go_in;
    logic tdcc_go_out;
    logic tdcc_done_in;
    logic tdcc_done_out;
    initial begin
        tcam_write_en = 1'd0;
        tcam_search_en = 1'd0;
        tcam_in = 32'd0;
        tcam_prefix_len = 6'd0;
        tcam_write_index = 5'd0;
        tcam_go = 1'd0;
        tcam_clk = 1'd0;
        tcam_reset = 1'd0;
        fsm_in = 2'd0;
        fsm_write_en = 1'd0;
        fsm_clk = 1'd0;
        fsm_reset = 1'd0;
        save_index_go_in = 1'd0;
        save_index_done_in = 1'd0;
        invoke_go_in = 1'd0;
        invoke_done_in = 1'd0;
        invoke0_go_in = 1'd0;
        invoke0_done_in = 1'd0;
        tdcc_go_in = 1'd0;
        tdcc_done_in = 1'd0;
    end
    TCAM_IPv4 tcam (
        .clk(tcam_clk),
        .done(tcam_done),
        .go(tcam_go),
        .in(tcam_in),
        .index(tcam_index),
        .prefix_len(tcam_prefix_len),
        .reset(tcam_reset),
        .search_en(tcam_search_en),
        .write_en(tcam_write_en),
        .write_index(tcam_write_index)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm (
        .clk(fsm_clk),
        .done(fsm_done),
        .in(fsm_in),
        .out(fsm_out),
        .reset(fsm_reset),
        .write_en(fsm_write_en)
    );
    std_wire # (
        .WIDTH(1)
    ) save_index_go (
        .in(save_index_go_in),
        .out(save_index_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) save_index_done (
        .in(save_index_done_in),
        .out(save_index_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke_go (
        .in(invoke_go_in),
        .out(invoke_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke_done (
        .in(invoke_done_in),
        .out(invoke_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke0_go (
        .in(invoke0_go_in),
        .out(invoke0_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke0_done (
        .in(invoke0_done_in),
        .out(invoke0_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc_go (
        .in(tdcc_go_in),
        .out(tdcc_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc_done (
        .in(tdcc_done_in),
        .out(tdcc_done_out)
    );
    assign done = tdcc_done_out;
    assign index_addr0 =
     save_index_go_out ? 1'd0 : 1'd0;
    assign index_clk = clk;
    assign index_write_data =
     save_index_go_out ? tcam_index : 5'd0;
    assign index_write_en = save_index_go_out;
    assign fsm_clk = clk;
    assign fsm_in =
     fsm_out == 2'd3 ? 2'd0 :
     fsm_out == 2'd0 & invoke_done_out & tdcc_go_out ? 2'd1 :
     fsm_out == 2'd1 & invoke0_done_out & tdcc_go_out ? 2'd2 :
     fsm_out == 2'd2 & save_index_done_out & tdcc_go_out ? 2'd3 : 2'd0;
    assign fsm_reset = reset;
    assign fsm_write_en = fsm_out == 2'd3 | fsm_out == 2'd0 & invoke_done_out & tdcc_go_out | fsm_out == 2'd1 & invoke0_done_out & tdcc_go_out | fsm_out == 2'd2 & save_index_done_out & tdcc_go_out;
    assign invoke0_done_in = tcam_done;
    assign invoke0_go_in = ~invoke0_done_out & fsm_out == 2'd1 & tdcc_go_out;
    assign invoke_done_in = tcam_done;
    assign invoke_go_in = ~invoke_done_out & fsm_out == 2'd0 & tdcc_go_out;
    assign save_index_done_in = index_done;
    assign save_index_go_in = ~save_index_done_out & fsm_out == 2'd2 & tdcc_go_out;
    assign tcam_clk = clk;
    assign tcam_go = invoke_go_out | invoke0_go_out;
    assign tcam_in =
     invoke_go_out ? 32'd0 :
     invoke0_go_out ? 32'd3221225472 : 32'd0;
    assign tcam_prefix_len =
     invoke_go_out ? 6'd0 : 6'd0;
    assign tcam_reset = reset;
    assign tcam_search_en = invoke0_go_out;
    assign tcam_write_en = invoke_go_out;
    assign tcam_write_index =
     invoke_go_out ? 5'd31 : 5'd0;
    assign tdcc_done_in = fsm_out == 2'd3;
    assign tdcc_go_in = go;
endmodule

module match_element (
    input logic [31:0] in,
    input logic [31:0] prefix,
    input logic [4:0] length,
    output logic out,
    input logic go,
    input logic clk,
    input logic reset,
    output logic done
);
    logic [4:0] sub_left;
    logic [4:0] sub_right;
    logic [4:0] sub_out;
    logic [4:0] pad_in;
    logic [31:0] pad_out;
    logic [31:0] rsh0_left;
    logic [31:0] rsh0_right;
    logic [31:0] rsh0_out;
    logic [31:0] rsh1_left;
    logic [31:0] rsh1_right;
    logic [31:0] rsh1_out;
    logic [31:0] eq_left;
    logic [31:0] eq_right;
    logic eq_out;
    logic r_in;
    logic r_write_en;
    logic r_clk;
    logic r_reset;
    logic r_out;
    logic r_done;
    logic compare_go_in;
    logic compare_go_out;
    logic compare_done_in;
    logic compare_done_out;
    initial begin
        sub_left = 5'd0;
        sub_right = 5'd0;
        pad_in = 5'd0;
        rsh0_left = 32'd0;
        rsh0_right = 32'd0;
        rsh1_left = 32'd0;
        rsh1_right = 32'd0;
        eq_left = 32'd0;
        eq_right = 32'd0;
        r_in = 1'd0;
        r_write_en = 1'd0;
        r_clk = 1'd0;
        r_reset = 1'd0;
        compare_go_in = 1'd0;
        compare_done_in = 1'd0;
    end
    std_sub # (
        .WIDTH(5)
    ) sub (
        .left(sub_left),
        .out(sub_out),
        .right(sub_right)
    );
    std_pad # (
        .IN_WIDTH(5),
        .OUT_WIDTH(32)
    ) pad (
        .in(pad_in),
        .out(pad_out)
    );
    std_rsh # (
        .WIDTH(32)
    ) rsh0 (
        .left(rsh0_left),
        .out(rsh0_out),
        .right(rsh0_right)
    );
    std_rsh # (
        .WIDTH(32)
    ) rsh1 (
        .left(rsh1_left),
        .out(rsh1_out),
        .right(rsh1_right)
    );
    std_eq # (
        .WIDTH(32)
    ) eq (
        .left(eq_left),
        .out(eq_out),
        .right(eq_right)
    );
    std_reg # (
        .WIDTH(1)
    ) r (
        .clk(r_clk),
        .done(r_done),
        .in(r_in),
        .out(r_out),
        .reset(r_reset),
        .write_en(r_write_en)
    );
    std_wire # (
        .WIDTH(1)
    ) compare_go (
        .in(compare_go_in),
        .out(compare_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) compare_done (
        .in(compare_done_in),
        .out(compare_done_out)
    );
    assign done = compare_done_out;
    assign out = r_out;
    assign compare_done_in = r_done;
    assign compare_go_in = go;
    assign eq_left =
     compare_go_out ? rsh0_out : 32'd0;
    assign eq_right =
     compare_go_out ? rsh1_out : 32'd0;
    assign pad_in =
     compare_go_out ? sub_out : 5'd0;
    assign r_clk = clk;
    assign r_in =
     compare_go_out ? eq_out : 1'd0;
    assign r_reset = reset;
    assign r_write_en = compare_go_out;
    assign rsh0_left =
     compare_go_out ? in : 32'd0;
    assign rsh0_right =
     compare_go_out ? pad_out : 32'd0;
    assign rsh1_left =
     compare_go_out ? prefix : 32'd0;
    assign rsh1_right =
     compare_go_out ? pad_out : 32'd0;
    assign sub_left =
     compare_go_out ? 5'd31 : 5'd0;
    assign sub_right =
     compare_go_out ? length : 5'd0;
endmodule

module comparator_element (
    input logic [4:0] lenA,
    input logic [4:0] lenB,
    input logic [4:0] addrA,
    input logic [4:0] addrB,
    input logic mlA,
    input logic mlB,
    output logic [4:0] lenX,
    output logic [4:0] addrX,
    output logic mlX,
    input logic go,
    input logic clk,
    input logic reset,
    output logic done
);
    logic [4:0] gt0_left;
    logic [4:0] gt0_right;
    logic gt0_out;
    logic or0_left;
    logic or0_right;
    logic or0_out;
    logic or1_left;
    logic or1_right;
    logic or1_out;
    logic not0_in;
    logic not0_out;
    logic and0_left;
    logic and0_right;
    logic and0_out;
    logic [4:0] len_in;
    logic len_write_en;
    logic len_clk;
    logic len_reset;
    logic [4:0] len_out;
    logic len_done;
    logic [4:0] addr_in;
    logic addr_write_en;
    logic addr_clk;
    logic addr_reset;
    logic [4:0] addr_out;
    logic addr_done;
    logic ml_in;
    logic ml_write_en;
    logic ml_clk;
    logic ml_reset;
    logic ml_out;
    logic ml_done;
    logic comb_reg_in;
    logic comb_reg_write_en;
    logic comb_reg_clk;
    logic comb_reg_reset;
    logic comb_reg_out;
    logic comb_reg_done;
    logic pd_in;
    logic pd_write_en;
    logic pd_clk;
    logic pd_reset;
    logic pd_out;
    logic pd_done;
    logic [1:0] fsm_in;
    logic fsm_write_en;
    logic fsm_clk;
    logic fsm_reset;
    logic [1:0] fsm_out;
    logic fsm_done;
    logic pd0_in;
    logic pd0_write_en;
    logic pd0_clk;
    logic pd0_reset;
    logic pd0_out;
    logic pd0_done;
    logic fsm0_in;
    logic fsm0_write_en;
    logic fsm0_clk;
    logic fsm0_reset;
    logic fsm0_out;
    logic fsm0_done;
    logic A_go_in;
    logic A_go_out;
    logic A_done_in;
    logic A_done_out;
    logic B_go_in;
    logic B_go_out;
    logic B_done_in;
    logic B_done_out;
    logic or_match_line_go_in;
    logic or_match_line_go_out;
    logic or_match_line_done_in;
    logic or_match_line_done_out;
    logic select0_go_in;
    logic select0_go_out;
    logic select0_done_in;
    logic select0_done_out;
    logic par_go_in;
    logic par_go_out;
    logic par_done_in;
    logic par_done_out;
    logic tdcc_go_in;
    logic tdcc_go_out;
    logic tdcc_done_in;
    logic tdcc_done_out;
    logic tdcc0_go_in;
    logic tdcc0_go_out;
    logic tdcc0_done_in;
    logic tdcc0_done_out;
    initial begin
        gt0_left = 5'd0;
        gt0_right = 5'd0;
        or0_left = 1'd0;
        or0_right = 1'd0;
        or1_left = 1'd0;
        or1_right = 1'd0;
        not0_in = 1'd0;
        and0_left = 1'd0;
        and0_right = 1'd0;
        len_in = 5'd0;
        len_write_en = 1'd0;
        len_clk = 1'd0;
        len_reset = 1'd0;
        addr_in = 5'd0;
        addr_write_en = 1'd0;
        addr_clk = 1'd0;
        addr_reset = 1'd0;
        ml_in = 1'd0;
        ml_write_en = 1'd0;
        ml_clk = 1'd0;
        ml_reset = 1'd0;
        comb_reg_in = 1'd0;
        comb_reg_write_en = 1'd0;
        comb_reg_clk = 1'd0;
        comb_reg_reset = 1'd0;
        pd_in = 1'd0;
        pd_write_en = 1'd0;
        pd_clk = 1'd0;
        pd_reset = 1'd0;
        fsm_in = 2'd0;
        fsm_write_en = 1'd0;
        fsm_clk = 1'd0;
        fsm_reset = 1'd0;
        pd0_in = 1'd0;
        pd0_write_en = 1'd0;
        pd0_clk = 1'd0;
        pd0_reset = 1'd0;
        fsm0_in = 1'd0;
        fsm0_write_en = 1'd0;
        fsm0_clk = 1'd0;
        fsm0_reset = 1'd0;
        A_go_in = 1'd0;
        A_done_in = 1'd0;
        B_go_in = 1'd0;
        B_done_in = 1'd0;
        or_match_line_go_in = 1'd0;
        or_match_line_done_in = 1'd0;
        select0_go_in = 1'd0;
        select0_done_in = 1'd0;
        par_go_in = 1'd0;
        par_done_in = 1'd0;
        tdcc_go_in = 1'd0;
        tdcc_done_in = 1'd0;
        tdcc0_go_in = 1'd0;
        tdcc0_done_in = 1'd0;
    end
    std_gt # (
        .WIDTH(5)
    ) gt0 (
        .left(gt0_left),
        .out(gt0_out),
        .right(gt0_right)
    );
    std_or # (
        .WIDTH(1)
    ) or0 (
        .left(or0_left),
        .out(or0_out),
        .right(or0_right)
    );
    std_or # (
        .WIDTH(1)
    ) or1 (
        .left(or1_left),
        .out(or1_out),
        .right(or1_right)
    );
    std_not # (
        .WIDTH(1)
    ) not0 (
        .in(not0_in),
        .out(not0_out)
    );
    std_and # (
        .WIDTH(1)
    ) and0 (
        .left(and0_left),
        .out(and0_out),
        .right(and0_right)
    );
    std_reg # (
        .WIDTH(5)
    ) len (
        .clk(len_clk),
        .done(len_done),
        .in(len_in),
        .out(len_out),
        .reset(len_reset),
        .write_en(len_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) addr (
        .clk(addr_clk),
        .done(addr_done),
        .in(addr_in),
        .out(addr_out),
        .reset(addr_reset),
        .write_en(addr_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) ml (
        .clk(ml_clk),
        .done(ml_done),
        .in(ml_in),
        .out(ml_out),
        .reset(ml_reset),
        .write_en(ml_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg (
        .clk(comb_reg_clk),
        .done(comb_reg_done),
        .in(comb_reg_in),
        .out(comb_reg_out),
        .reset(comb_reg_reset),
        .write_en(comb_reg_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd (
        .clk(pd_clk),
        .done(pd_done),
        .in(pd_in),
        .out(pd_out),
        .reset(pd_reset),
        .write_en(pd_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm (
        .clk(fsm_clk),
        .done(fsm_done),
        .in(fsm_in),
        .out(fsm_out),
        .reset(fsm_reset),
        .write_en(fsm_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd0 (
        .clk(pd0_clk),
        .done(pd0_done),
        .in(pd0_in),
        .out(pd0_out),
        .reset(pd0_reset),
        .write_en(pd0_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) fsm0 (
        .clk(fsm0_clk),
        .done(fsm0_done),
        .in(fsm0_in),
        .out(fsm0_out),
        .reset(fsm0_reset),
        .write_en(fsm0_write_en)
    );
    std_wire # (
        .WIDTH(1)
    ) A_go (
        .in(A_go_in),
        .out(A_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) A_done (
        .in(A_done_in),
        .out(A_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) B_go (
        .in(B_go_in),
        .out(B_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) B_done (
        .in(B_done_in),
        .out(B_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) or_match_line_go (
        .in(or_match_line_go_in),
        .out(or_match_line_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) or_match_line_done (
        .in(or_match_line_done_in),
        .out(or_match_line_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) select0_go (
        .in(select0_go_in),
        .out(select0_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) select0_done (
        .in(select0_done_in),
        .out(select0_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par_go (
        .in(par_go_in),
        .out(par_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par_done (
        .in(par_done_in),
        .out(par_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc_go (
        .in(tdcc_go_in),
        .out(tdcc_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc_done (
        .in(tdcc_done_in),
        .out(tdcc_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc0_go (
        .in(tdcc0_go_in),
        .out(tdcc0_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc0_done (
        .in(tdcc0_done_in),
        .out(tdcc0_done_out)
    );
    assign A_done_in = len_done & addr_done;
    assign A_go_in = ~A_done_out & fsm_out == 2'd1 & tdcc_go_out;
    assign B_done_in = len_done & addr_done;
    assign B_go_in = ~B_done_out & fsm_out == 2'd2 & tdcc_go_out;
    assign addrX = addr_out;
    assign done = tdcc0_done_out;
    assign lenX = len_out;
    assign mlX = ml_out;
    assign addr_clk = clk;
    assign addr_in =
     A_go_out ? addrA :
     B_go_out ? addrB : 5'd0;
    assign addr_reset = reset;
    assign addr_write_en = A_go_out | B_go_out;
    assign and0_left =
     select0_go_out ? mlA : 1'd0;
    assign and0_right =
     select0_go_out ? or0_out : 1'd0;
    assign comb_reg_clk = clk;
    assign comb_reg_in =
     select0_go_out ? and0_out : 1'd0;
    assign comb_reg_reset = reset;
    assign comb_reg_write_en = select0_go_out;
    assign fsm_clk = clk;
    assign fsm_in =
     fsm_out == 2'd3 ? 2'd0 :
     fsm_out == 2'd0 & select0_done_out & comb_reg_out & tdcc_go_out ? 2'd1 :
     fsm_out == 2'd0 & select0_done_out & ~comb_reg_out & tdcc_go_out ? 2'd2 :
     fsm_out == 2'd1 & A_done_out & tdcc_go_out | fsm_out == 2'd2 & B_done_out & tdcc_go_out ? 2'd3 : 2'd0;
    assign fsm_reset = reset;
    assign fsm_write_en = fsm_out == 2'd3 | fsm_out == 2'd0 & select0_done_out & comb_reg_out & tdcc_go_out | fsm_out == 2'd0 & select0_done_out & ~comb_reg_out & tdcc_go_out | fsm_out == 2'd1 & A_done_out & tdcc_go_out | fsm_out == 2'd2 & B_done_out & tdcc_go_out;
    assign fsm0_clk = clk;
    assign fsm0_in =
     fsm0_out == 1'd1 ? 1'd0 :
     fsm0_out == 1'd0 & par_done_out & tdcc0_go_out ? 1'd1 : 1'd0;
    assign fsm0_reset = reset;
    assign fsm0_write_en = fsm0_out == 1'd1 | fsm0_out == 1'd0 & par_done_out & tdcc0_go_out;
    assign gt0_left =
     select0_go_out ? lenA : 5'd0;
    assign gt0_right =
     select0_go_out ? lenB : 5'd0;
    assign len_clk = clk;
    assign len_in =
     A_go_out ? lenA :
     B_go_out ? lenB : 5'd0;
    assign len_reset = reset;
    assign len_write_en = A_go_out | B_go_out;
    assign ml_clk = clk;
    assign ml_in =
     or_match_line_go_out ? or1_out : 1'd0;
    assign ml_reset = reset;
    assign ml_write_en = or_match_line_go_out;
    assign not0_in =
     select0_go_out ? mlB : 1'd0;
    assign or0_left =
     select0_go_out ? not0_out : 1'd0;
    assign or0_right =
     select0_go_out ? gt0_out : 1'd0;
    assign or1_left =
     or_match_line_go_out ? mlA : 1'd0;
    assign or1_right =
     or_match_line_go_out ? mlB : 1'd0;
    assign or_match_line_done_in = ml_done;
    assign or_match_line_go_in = ~(pd_out | or_match_line_done_out) & par_go_out;
    assign par_done_in = pd_out & pd0_out;
    assign par_go_in = ~par_done_out & fsm0_out == 1'd0 & tdcc0_go_out;
    assign pd_clk = clk;
    assign pd_in =
     pd_out & pd0_out ? 1'd0 :
     or_match_line_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd_reset = reset;
    assign pd_write_en = pd_out & pd0_out | or_match_line_done_out & par_go_out;
    assign pd0_clk = clk;
    assign pd0_in =
     pd_out & pd0_out ? 1'd0 :
     tdcc_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd0_reset = reset;
    assign pd0_write_en = pd_out & pd0_out | tdcc_done_out & par_go_out;
    assign select0_done_in = comb_reg_done;
    assign select0_go_in = ~select0_done_out & fsm_out == 2'd0 & tdcc_go_out;
    assign tdcc0_done_in = fsm0_out == 1'd1;
    assign tdcc0_go_in = go;
    assign tdcc_done_in = fsm_out == 2'd3;
    assign tdcc_go_in = ~(pd0_out | tdcc_done_out) & par_go_out;
endmodule

module TCAM_IPv4 (
    input logic write_en,
    input logic search_en,
    input logic [31:0] in,
    input logic [5:0] prefix_len,
    input logic [4:0] write_index,
    output logic [4:0] index,
    input logic go,
    input logic clk,
    input logic reset,
    output logic done
);
    logic [31:0] p0_in;
    logic p0_write_en;
    logic p0_clk;
    logic p0_reset;
    logic [31:0] p0_out;
    logic p0_done;
    logic [31:0] p1_in;
    logic p1_write_en;
    logic p1_clk;
    logic p1_reset;
    logic [31:0] p1_out;
    logic p1_done;
    logic [31:0] p2_in;
    logic p2_write_en;
    logic p2_clk;
    logic p2_reset;
    logic [31:0] p2_out;
    logic p2_done;
    logic [31:0] p3_in;
    logic p3_write_en;
    logic p3_clk;
    logic p3_reset;
    logic [31:0] p3_out;
    logic p3_done;
    logic [31:0] p4_in;
    logic p4_write_en;
    logic p4_clk;
    logic p4_reset;
    logic [31:0] p4_out;
    logic p4_done;
    logic [31:0] p5_in;
    logic p5_write_en;
    logic p5_clk;
    logic p5_reset;
    logic [31:0] p5_out;
    logic p5_done;
    logic [31:0] p6_in;
    logic p6_write_en;
    logic p6_clk;
    logic p6_reset;
    logic [31:0] p6_out;
    logic p6_done;
    logic [31:0] p7_in;
    logic p7_write_en;
    logic p7_clk;
    logic p7_reset;
    logic [31:0] p7_out;
    logic p7_done;
    logic [31:0] p8_in;
    logic p8_write_en;
    logic p8_clk;
    logic p8_reset;
    logic [31:0] p8_out;
    logic p8_done;
    logic [31:0] p9_in;
    logic p9_write_en;
    logic p9_clk;
    logic p9_reset;
    logic [31:0] p9_out;
    logic p9_done;
    logic [31:0] p10_in;
    logic p10_write_en;
    logic p10_clk;
    logic p10_reset;
    logic [31:0] p10_out;
    logic p10_done;
    logic [31:0] p11_in;
    logic p11_write_en;
    logic p11_clk;
    logic p11_reset;
    logic [31:0] p11_out;
    logic p11_done;
    logic [31:0] p12_in;
    logic p12_write_en;
    logic p12_clk;
    logic p12_reset;
    logic [31:0] p12_out;
    logic p12_done;
    logic [31:0] p13_in;
    logic p13_write_en;
    logic p13_clk;
    logic p13_reset;
    logic [31:0] p13_out;
    logic p13_done;
    logic [31:0] p14_in;
    logic p14_write_en;
    logic p14_clk;
    logic p14_reset;
    logic [31:0] p14_out;
    logic p14_done;
    logic [31:0] p15_in;
    logic p15_write_en;
    logic p15_clk;
    logic p15_reset;
    logic [31:0] p15_out;
    logic p15_done;
    logic [31:0] p16_in;
    logic p16_write_en;
    logic p16_clk;
    logic p16_reset;
    logic [31:0] p16_out;
    logic p16_done;
    logic [31:0] p17_in;
    logic p17_write_en;
    logic p17_clk;
    logic p17_reset;
    logic [31:0] p17_out;
    logic p17_done;
    logic [31:0] p18_in;
    logic p18_write_en;
    logic p18_clk;
    logic p18_reset;
    logic [31:0] p18_out;
    logic p18_done;
    logic [31:0] p19_in;
    logic p19_write_en;
    logic p19_clk;
    logic p19_reset;
    logic [31:0] p19_out;
    logic p19_done;
    logic [31:0] p20_in;
    logic p20_write_en;
    logic p20_clk;
    logic p20_reset;
    logic [31:0] p20_out;
    logic p20_done;
    logic [31:0] p21_in;
    logic p21_write_en;
    logic p21_clk;
    logic p21_reset;
    logic [31:0] p21_out;
    logic p21_done;
    logic [31:0] p22_in;
    logic p22_write_en;
    logic p22_clk;
    logic p22_reset;
    logic [31:0] p22_out;
    logic p22_done;
    logic [31:0] p23_in;
    logic p23_write_en;
    logic p23_clk;
    logic p23_reset;
    logic [31:0] p23_out;
    logic p23_done;
    logic [31:0] p24_in;
    logic p24_write_en;
    logic p24_clk;
    logic p24_reset;
    logic [31:0] p24_out;
    logic p24_done;
    logic [31:0] p25_in;
    logic p25_write_en;
    logic p25_clk;
    logic p25_reset;
    logic [31:0] p25_out;
    logic p25_done;
    logic [31:0] p26_in;
    logic p26_write_en;
    logic p26_clk;
    logic p26_reset;
    logic [31:0] p26_out;
    logic p26_done;
    logic [31:0] p27_in;
    logic p27_write_en;
    logic p27_clk;
    logic p27_reset;
    logic [31:0] p27_out;
    logic p27_done;
    logic [31:0] p28_in;
    logic p28_write_en;
    logic p28_clk;
    logic p28_reset;
    logic [31:0] p28_out;
    logic p28_done;
    logic [31:0] p29_in;
    logic p29_write_en;
    logic p29_clk;
    logic p29_reset;
    logic [31:0] p29_out;
    logic p29_done;
    logic [31:0] p30_in;
    logic p30_write_en;
    logic p30_clk;
    logic p30_reset;
    logic [31:0] p30_out;
    logic p30_done;
    logic [31:0] p31_in;
    logic p31_write_en;
    logic p31_clk;
    logic p31_reset;
    logic [31:0] p31_out;
    logic p31_done;
    logic [4:0] l0_in;
    logic l0_write_en;
    logic l0_clk;
    logic l0_reset;
    logic [4:0] l0_out;
    logic l0_done;
    logic [4:0] l1_in;
    logic l1_write_en;
    logic l1_clk;
    logic l1_reset;
    logic [4:0] l1_out;
    logic l1_done;
    logic [4:0] l2_in;
    logic l2_write_en;
    logic l2_clk;
    logic l2_reset;
    logic [4:0] l2_out;
    logic l2_done;
    logic [4:0] l3_in;
    logic l3_write_en;
    logic l3_clk;
    logic l3_reset;
    logic [4:0] l3_out;
    logic l3_done;
    logic [4:0] l4_in;
    logic l4_write_en;
    logic l4_clk;
    logic l4_reset;
    logic [4:0] l4_out;
    logic l4_done;
    logic [4:0] l5_in;
    logic l5_write_en;
    logic l5_clk;
    logic l5_reset;
    logic [4:0] l5_out;
    logic l5_done;
    logic [4:0] l6_in;
    logic l6_write_en;
    logic l6_clk;
    logic l6_reset;
    logic [4:0] l6_out;
    logic l6_done;
    logic [4:0] l7_in;
    logic l7_write_en;
    logic l7_clk;
    logic l7_reset;
    logic [4:0] l7_out;
    logic l7_done;
    logic [4:0] l8_in;
    logic l8_write_en;
    logic l8_clk;
    logic l8_reset;
    logic [4:0] l8_out;
    logic l8_done;
    logic [4:0] l9_in;
    logic l9_write_en;
    logic l9_clk;
    logic l9_reset;
    logic [4:0] l9_out;
    logic l9_done;
    logic [4:0] l10_in;
    logic l10_write_en;
    logic l10_clk;
    logic l10_reset;
    logic [4:0] l10_out;
    logic l10_done;
    logic [4:0] l11_in;
    logic l11_write_en;
    logic l11_clk;
    logic l11_reset;
    logic [4:0] l11_out;
    logic l11_done;
    logic [4:0] l12_in;
    logic l12_write_en;
    logic l12_clk;
    logic l12_reset;
    logic [4:0] l12_out;
    logic l12_done;
    logic [4:0] l13_in;
    logic l13_write_en;
    logic l13_clk;
    logic l13_reset;
    logic [4:0] l13_out;
    logic l13_done;
    logic [4:0] l14_in;
    logic l14_write_en;
    logic l14_clk;
    logic l14_reset;
    logic [4:0] l14_out;
    logic l14_done;
    logic [4:0] l15_in;
    logic l15_write_en;
    logic l15_clk;
    logic l15_reset;
    logic [4:0] l15_out;
    logic l15_done;
    logic [4:0] l16_in;
    logic l16_write_en;
    logic l16_clk;
    logic l16_reset;
    logic [4:0] l16_out;
    logic l16_done;
    logic [4:0] l17_in;
    logic l17_write_en;
    logic l17_clk;
    logic l17_reset;
    logic [4:0] l17_out;
    logic l17_done;
    logic [4:0] l18_in;
    logic l18_write_en;
    logic l18_clk;
    logic l18_reset;
    logic [4:0] l18_out;
    logic l18_done;
    logic [4:0] l19_in;
    logic l19_write_en;
    logic l19_clk;
    logic l19_reset;
    logic [4:0] l19_out;
    logic l19_done;
    logic [4:0] l20_in;
    logic l20_write_en;
    logic l20_clk;
    logic l20_reset;
    logic [4:0] l20_out;
    logic l20_done;
    logic [4:0] l21_in;
    logic l21_write_en;
    logic l21_clk;
    logic l21_reset;
    logic [4:0] l21_out;
    logic l21_done;
    logic [4:0] l22_in;
    logic l22_write_en;
    logic l22_clk;
    logic l22_reset;
    logic [4:0] l22_out;
    logic l22_done;
    logic [4:0] l23_in;
    logic l23_write_en;
    logic l23_clk;
    logic l23_reset;
    logic [4:0] l23_out;
    logic l23_done;
    logic [4:0] l24_in;
    logic l24_write_en;
    logic l24_clk;
    logic l24_reset;
    logic [4:0] l24_out;
    logic l24_done;
    logic [4:0] l25_in;
    logic l25_write_en;
    logic l25_clk;
    logic l25_reset;
    logic [4:0] l25_out;
    logic l25_done;
    logic [4:0] l26_in;
    logic l26_write_en;
    logic l26_clk;
    logic l26_reset;
    logic [4:0] l26_out;
    logic l26_done;
    logic [4:0] l27_in;
    logic l27_write_en;
    logic l27_clk;
    logic l27_reset;
    logic [4:0] l27_out;
    logic l27_done;
    logic [4:0] l28_in;
    logic l28_write_en;
    logic l28_clk;
    logic l28_reset;
    logic [4:0] l28_out;
    logic l28_done;
    logic [4:0] l29_in;
    logic l29_write_en;
    logic l29_clk;
    logic l29_reset;
    logic [4:0] l29_out;
    logic l29_done;
    logic [4:0] l30_in;
    logic l30_write_en;
    logic l30_clk;
    logic l30_reset;
    logic [4:0] l30_out;
    logic l30_done;
    logic [4:0] l31_in;
    logic l31_write_en;
    logic l31_clk;
    logic l31_reset;
    logic [4:0] l31_out;
    logic l31_done;
    logic [4:0] is_index0_left;
    logic [4:0] is_index0_right;
    logic is_index0_out;
    logic [4:0] is_index1_left;
    logic [4:0] is_index1_right;
    logic is_index1_out;
    logic [4:0] is_index2_left;
    logic [4:0] is_index2_right;
    logic is_index2_out;
    logic [4:0] is_index3_left;
    logic [4:0] is_index3_right;
    logic is_index3_out;
    logic [4:0] is_index4_left;
    logic [4:0] is_index4_right;
    logic is_index4_out;
    logic [4:0] is_index5_left;
    logic [4:0] is_index5_right;
    logic is_index5_out;
    logic [4:0] is_index6_left;
    logic [4:0] is_index6_right;
    logic is_index6_out;
    logic [4:0] is_index7_left;
    logic [4:0] is_index7_right;
    logic is_index7_out;
    logic [4:0] is_index8_left;
    logic [4:0] is_index8_right;
    logic is_index8_out;
    logic [4:0] is_index9_left;
    logic [4:0] is_index9_right;
    logic is_index9_out;
    logic [4:0] is_index10_left;
    logic [4:0] is_index10_right;
    logic is_index10_out;
    logic [4:0] is_index11_left;
    logic [4:0] is_index11_right;
    logic is_index11_out;
    logic [4:0] is_index12_left;
    logic [4:0] is_index12_right;
    logic is_index12_out;
    logic [4:0] is_index13_left;
    logic [4:0] is_index13_right;
    logic is_index13_out;
    logic [4:0] is_index14_left;
    logic [4:0] is_index14_right;
    logic is_index14_out;
    logic [4:0] is_index15_left;
    logic [4:0] is_index15_right;
    logic is_index15_out;
    logic [4:0] is_index16_left;
    logic [4:0] is_index16_right;
    logic is_index16_out;
    logic [4:0] is_index17_left;
    logic [4:0] is_index17_right;
    logic is_index17_out;
    logic [4:0] is_index18_left;
    logic [4:0] is_index18_right;
    logic is_index18_out;
    logic [4:0] is_index19_left;
    logic [4:0] is_index19_right;
    logic is_index19_out;
    logic [4:0] is_index20_left;
    logic [4:0] is_index20_right;
    logic is_index20_out;
    logic [4:0] is_index21_left;
    logic [4:0] is_index21_right;
    logic is_index21_out;
    logic [4:0] is_index22_left;
    logic [4:0] is_index22_right;
    logic is_index22_out;
    logic [4:0] is_index23_left;
    logic [4:0] is_index23_right;
    logic is_index23_out;
    logic [4:0] is_index24_left;
    logic [4:0] is_index24_right;
    logic is_index24_out;
    logic [4:0] is_index25_left;
    logic [4:0] is_index25_right;
    logic is_index25_out;
    logic [4:0] is_index26_left;
    logic [4:0] is_index26_right;
    logic is_index26_out;
    logic [4:0] is_index27_left;
    logic [4:0] is_index27_right;
    logic is_index27_out;
    logic [4:0] is_index28_left;
    logic [4:0] is_index28_right;
    logic is_index28_out;
    logic [4:0] is_index29_left;
    logic [4:0] is_index29_right;
    logic is_index29_out;
    logic [4:0] is_index30_left;
    logic [4:0] is_index30_right;
    logic is_index30_out;
    logic [4:0] is_index31_left;
    logic [4:0] is_index31_right;
    logic is_index31_out;
    logic [4:0] zero_index_in;
    logic zero_index_write_en;
    logic zero_index_clk;
    logic zero_index_reset;
    logic [4:0] zero_index_out;
    logic zero_index_done;
    logic [5:0] z_eq_left;
    logic [5:0] z_eq_right;
    logic z_eq_out;
    logic [5:0] slice_in;
    logic [4:0] slice_out;
    logic [5:0] sub_left;
    logic [5:0] sub_right;
    logic [5:0] sub_out;
    logic [31:0] me0_in;
    logic [31:0] me0_prefix;
    logic [4:0] me0_length;
    logic me0_out;
    logic me0_go;
    logic me0_clk;
    logic me0_reset;
    logic me0_done;
    logic [31:0] me1_in;
    logic [31:0] me1_prefix;
    logic [4:0] me1_length;
    logic me1_out;
    logic me1_go;
    logic me1_clk;
    logic me1_reset;
    logic me1_done;
    logic [31:0] me2_in;
    logic [31:0] me2_prefix;
    logic [4:0] me2_length;
    logic me2_out;
    logic me2_go;
    logic me2_clk;
    logic me2_reset;
    logic me2_done;
    logic [31:0] me3_in;
    logic [31:0] me3_prefix;
    logic [4:0] me3_length;
    logic me3_out;
    logic me3_go;
    logic me3_clk;
    logic me3_reset;
    logic me3_done;
    logic [31:0] me4_in;
    logic [31:0] me4_prefix;
    logic [4:0] me4_length;
    logic me4_out;
    logic me4_go;
    logic me4_clk;
    logic me4_reset;
    logic me4_done;
    logic [31:0] me5_in;
    logic [31:0] me5_prefix;
    logic [4:0] me5_length;
    logic me5_out;
    logic me5_go;
    logic me5_clk;
    logic me5_reset;
    logic me5_done;
    logic [31:0] me6_in;
    logic [31:0] me6_prefix;
    logic [4:0] me6_length;
    logic me6_out;
    logic me6_go;
    logic me6_clk;
    logic me6_reset;
    logic me6_done;
    logic [31:0] me7_in;
    logic [31:0] me7_prefix;
    logic [4:0] me7_length;
    logic me7_out;
    logic me7_go;
    logic me7_clk;
    logic me7_reset;
    logic me7_done;
    logic [31:0] me8_in;
    logic [31:0] me8_prefix;
    logic [4:0] me8_length;
    logic me8_out;
    logic me8_go;
    logic me8_clk;
    logic me8_reset;
    logic me8_done;
    logic [31:0] me9_in;
    logic [31:0] me9_prefix;
    logic [4:0] me9_length;
    logic me9_out;
    logic me9_go;
    logic me9_clk;
    logic me9_reset;
    logic me9_done;
    logic [31:0] me10_in;
    logic [31:0] me10_prefix;
    logic [4:0] me10_length;
    logic me10_out;
    logic me10_go;
    logic me10_clk;
    logic me10_reset;
    logic me10_done;
    logic [31:0] me11_in;
    logic [31:0] me11_prefix;
    logic [4:0] me11_length;
    logic me11_out;
    logic me11_go;
    logic me11_clk;
    logic me11_reset;
    logic me11_done;
    logic [31:0] me12_in;
    logic [31:0] me12_prefix;
    logic [4:0] me12_length;
    logic me12_out;
    logic me12_go;
    logic me12_clk;
    logic me12_reset;
    logic me12_done;
    logic [31:0] me13_in;
    logic [31:0] me13_prefix;
    logic [4:0] me13_length;
    logic me13_out;
    logic me13_go;
    logic me13_clk;
    logic me13_reset;
    logic me13_done;
    logic [31:0] me14_in;
    logic [31:0] me14_prefix;
    logic [4:0] me14_length;
    logic me14_out;
    logic me14_go;
    logic me14_clk;
    logic me14_reset;
    logic me14_done;
    logic [31:0] me15_in;
    logic [31:0] me15_prefix;
    logic [4:0] me15_length;
    logic me15_out;
    logic me15_go;
    logic me15_clk;
    logic me15_reset;
    logic me15_done;
    logic [31:0] me16_in;
    logic [31:0] me16_prefix;
    logic [4:0] me16_length;
    logic me16_out;
    logic me16_go;
    logic me16_clk;
    logic me16_reset;
    logic me16_done;
    logic [31:0] me17_in;
    logic [31:0] me17_prefix;
    logic [4:0] me17_length;
    logic me17_out;
    logic me17_go;
    logic me17_clk;
    logic me17_reset;
    logic me17_done;
    logic [31:0] me18_in;
    logic [31:0] me18_prefix;
    logic [4:0] me18_length;
    logic me18_out;
    logic me18_go;
    logic me18_clk;
    logic me18_reset;
    logic me18_done;
    logic [31:0] me19_in;
    logic [31:0] me19_prefix;
    logic [4:0] me19_length;
    logic me19_out;
    logic me19_go;
    logic me19_clk;
    logic me19_reset;
    logic me19_done;
    logic [31:0] me20_in;
    logic [31:0] me20_prefix;
    logic [4:0] me20_length;
    logic me20_out;
    logic me20_go;
    logic me20_clk;
    logic me20_reset;
    logic me20_done;
    logic [31:0] me21_in;
    logic [31:0] me21_prefix;
    logic [4:0] me21_length;
    logic me21_out;
    logic me21_go;
    logic me21_clk;
    logic me21_reset;
    logic me21_done;
    logic [31:0] me22_in;
    logic [31:0] me22_prefix;
    logic [4:0] me22_length;
    logic me22_out;
    logic me22_go;
    logic me22_clk;
    logic me22_reset;
    logic me22_done;
    logic [31:0] me23_in;
    logic [31:0] me23_prefix;
    logic [4:0] me23_length;
    logic me23_out;
    logic me23_go;
    logic me23_clk;
    logic me23_reset;
    logic me23_done;
    logic [31:0] me24_in;
    logic [31:0] me24_prefix;
    logic [4:0] me24_length;
    logic me24_out;
    logic me24_go;
    logic me24_clk;
    logic me24_reset;
    logic me24_done;
    logic [31:0] me25_in;
    logic [31:0] me25_prefix;
    logic [4:0] me25_length;
    logic me25_out;
    logic me25_go;
    logic me25_clk;
    logic me25_reset;
    logic me25_done;
    logic [31:0] me26_in;
    logic [31:0] me26_prefix;
    logic [4:0] me26_length;
    logic me26_out;
    logic me26_go;
    logic me26_clk;
    logic me26_reset;
    logic me26_done;
    logic [31:0] me27_in;
    logic [31:0] me27_prefix;
    logic [4:0] me27_length;
    logic me27_out;
    logic me27_go;
    logic me27_clk;
    logic me27_reset;
    logic me27_done;
    logic [31:0] me28_in;
    logic [31:0] me28_prefix;
    logic [4:0] me28_length;
    logic me28_out;
    logic me28_go;
    logic me28_clk;
    logic me28_reset;
    logic me28_done;
    logic [31:0] me29_in;
    logic [31:0] me29_prefix;
    logic [4:0] me29_length;
    logic me29_out;
    logic me29_go;
    logic me29_clk;
    logic me29_reset;
    logic me29_done;
    logic [31:0] me30_in;
    logic [31:0] me30_prefix;
    logic [4:0] me30_length;
    logic me30_out;
    logic me30_go;
    logic me30_clk;
    logic me30_reset;
    logic me30_done;
    logic [31:0] me31_in;
    logic [31:0] me31_prefix;
    logic [4:0] me31_length;
    logic me31_out;
    logic me31_go;
    logic me31_clk;
    logic me31_reset;
    logic me31_done;
    logic [4:0] ce00_lenA;
    logic [4:0] ce00_lenB;
    logic [4:0] ce00_addrA;
    logic [4:0] ce00_addrB;
    logic ce00_mlA;
    logic ce00_mlB;
    logic [4:0] ce00_lenX;
    logic [4:0] ce00_addrX;
    logic ce00_mlX;
    logic ce00_go;
    logic ce00_clk;
    logic ce00_reset;
    logic ce00_done;
    logic [4:0] ce01_lenA;
    logic [4:0] ce01_lenB;
    logic [4:0] ce01_addrA;
    logic [4:0] ce01_addrB;
    logic ce01_mlA;
    logic ce01_mlB;
    logic [4:0] ce01_lenX;
    logic [4:0] ce01_addrX;
    logic ce01_mlX;
    logic ce01_go;
    logic ce01_clk;
    logic ce01_reset;
    logic ce01_done;
    logic [4:0] ce02_lenA;
    logic [4:0] ce02_lenB;
    logic [4:0] ce02_addrA;
    logic [4:0] ce02_addrB;
    logic ce02_mlA;
    logic ce02_mlB;
    logic [4:0] ce02_lenX;
    logic [4:0] ce02_addrX;
    logic ce02_mlX;
    logic ce02_go;
    logic ce02_clk;
    logic ce02_reset;
    logic ce02_done;
    logic [4:0] ce03_lenA;
    logic [4:0] ce03_lenB;
    logic [4:0] ce03_addrA;
    logic [4:0] ce03_addrB;
    logic ce03_mlA;
    logic ce03_mlB;
    logic [4:0] ce03_lenX;
    logic [4:0] ce03_addrX;
    logic ce03_mlX;
    logic ce03_go;
    logic ce03_clk;
    logic ce03_reset;
    logic ce03_done;
    logic [4:0] ce04_lenA;
    logic [4:0] ce04_lenB;
    logic [4:0] ce04_addrA;
    logic [4:0] ce04_addrB;
    logic ce04_mlA;
    logic ce04_mlB;
    logic [4:0] ce04_lenX;
    logic [4:0] ce04_addrX;
    logic ce04_mlX;
    logic ce04_go;
    logic ce04_clk;
    logic ce04_reset;
    logic ce04_done;
    logic [4:0] ce05_lenA;
    logic [4:0] ce05_lenB;
    logic [4:0] ce05_addrA;
    logic [4:0] ce05_addrB;
    logic ce05_mlA;
    logic ce05_mlB;
    logic [4:0] ce05_lenX;
    logic [4:0] ce05_addrX;
    logic ce05_mlX;
    logic ce05_go;
    logic ce05_clk;
    logic ce05_reset;
    logic ce05_done;
    logic [4:0] ce06_lenA;
    logic [4:0] ce06_lenB;
    logic [4:0] ce06_addrA;
    logic [4:0] ce06_addrB;
    logic ce06_mlA;
    logic ce06_mlB;
    logic [4:0] ce06_lenX;
    logic [4:0] ce06_addrX;
    logic ce06_mlX;
    logic ce06_go;
    logic ce06_clk;
    logic ce06_reset;
    logic ce06_done;
    logic [4:0] ce07_lenA;
    logic [4:0] ce07_lenB;
    logic [4:0] ce07_addrA;
    logic [4:0] ce07_addrB;
    logic ce07_mlA;
    logic ce07_mlB;
    logic [4:0] ce07_lenX;
    logic [4:0] ce07_addrX;
    logic ce07_mlX;
    logic ce07_go;
    logic ce07_clk;
    logic ce07_reset;
    logic ce07_done;
    logic [4:0] ce08_lenA;
    logic [4:0] ce08_lenB;
    logic [4:0] ce08_addrA;
    logic [4:0] ce08_addrB;
    logic ce08_mlA;
    logic ce08_mlB;
    logic [4:0] ce08_lenX;
    logic [4:0] ce08_addrX;
    logic ce08_mlX;
    logic ce08_go;
    logic ce08_clk;
    logic ce08_reset;
    logic ce08_done;
    logic [4:0] ce09_lenA;
    logic [4:0] ce09_lenB;
    logic [4:0] ce09_addrA;
    logic [4:0] ce09_addrB;
    logic ce09_mlA;
    logic ce09_mlB;
    logic [4:0] ce09_lenX;
    logic [4:0] ce09_addrX;
    logic ce09_mlX;
    logic ce09_go;
    logic ce09_clk;
    logic ce09_reset;
    logic ce09_done;
    logic [4:0] ce010_lenA;
    logic [4:0] ce010_lenB;
    logic [4:0] ce010_addrA;
    logic [4:0] ce010_addrB;
    logic ce010_mlA;
    logic ce010_mlB;
    logic [4:0] ce010_lenX;
    logic [4:0] ce010_addrX;
    logic ce010_mlX;
    logic ce010_go;
    logic ce010_clk;
    logic ce010_reset;
    logic ce010_done;
    logic [4:0] ce011_lenA;
    logic [4:0] ce011_lenB;
    logic [4:0] ce011_addrA;
    logic [4:0] ce011_addrB;
    logic ce011_mlA;
    logic ce011_mlB;
    logic [4:0] ce011_lenX;
    logic [4:0] ce011_addrX;
    logic ce011_mlX;
    logic ce011_go;
    logic ce011_clk;
    logic ce011_reset;
    logic ce011_done;
    logic [4:0] ce012_lenA;
    logic [4:0] ce012_lenB;
    logic [4:0] ce012_addrA;
    logic [4:0] ce012_addrB;
    logic ce012_mlA;
    logic ce012_mlB;
    logic [4:0] ce012_lenX;
    logic [4:0] ce012_addrX;
    logic ce012_mlX;
    logic ce012_go;
    logic ce012_clk;
    logic ce012_reset;
    logic ce012_done;
    logic [4:0] ce013_lenA;
    logic [4:0] ce013_lenB;
    logic [4:0] ce013_addrA;
    logic [4:0] ce013_addrB;
    logic ce013_mlA;
    logic ce013_mlB;
    logic [4:0] ce013_lenX;
    logic [4:0] ce013_addrX;
    logic ce013_mlX;
    logic ce013_go;
    logic ce013_clk;
    logic ce013_reset;
    logic ce013_done;
    logic [4:0] ce014_lenA;
    logic [4:0] ce014_lenB;
    logic [4:0] ce014_addrA;
    logic [4:0] ce014_addrB;
    logic ce014_mlA;
    logic ce014_mlB;
    logic [4:0] ce014_lenX;
    logic [4:0] ce014_addrX;
    logic ce014_mlX;
    logic ce014_go;
    logic ce014_clk;
    logic ce014_reset;
    logic ce014_done;
    logic [4:0] ce015_lenA;
    logic [4:0] ce015_lenB;
    logic [4:0] ce015_addrA;
    logic [4:0] ce015_addrB;
    logic ce015_mlA;
    logic ce015_mlB;
    logic [4:0] ce015_lenX;
    logic [4:0] ce015_addrX;
    logic ce015_mlX;
    logic ce015_go;
    logic ce015_clk;
    logic ce015_reset;
    logic ce015_done;
    logic [4:0] ce10_lenA;
    logic [4:0] ce10_lenB;
    logic [4:0] ce10_addrA;
    logic [4:0] ce10_addrB;
    logic ce10_mlA;
    logic ce10_mlB;
    logic [4:0] ce10_lenX;
    logic [4:0] ce10_addrX;
    logic ce10_mlX;
    logic ce10_go;
    logic ce10_clk;
    logic ce10_reset;
    logic ce10_done;
    logic [4:0] ce11_lenA;
    logic [4:0] ce11_lenB;
    logic [4:0] ce11_addrA;
    logic [4:0] ce11_addrB;
    logic ce11_mlA;
    logic ce11_mlB;
    logic [4:0] ce11_lenX;
    logic [4:0] ce11_addrX;
    logic ce11_mlX;
    logic ce11_go;
    logic ce11_clk;
    logic ce11_reset;
    logic ce11_done;
    logic [4:0] ce12_lenA;
    logic [4:0] ce12_lenB;
    logic [4:0] ce12_addrA;
    logic [4:0] ce12_addrB;
    logic ce12_mlA;
    logic ce12_mlB;
    logic [4:0] ce12_lenX;
    logic [4:0] ce12_addrX;
    logic ce12_mlX;
    logic ce12_go;
    logic ce12_clk;
    logic ce12_reset;
    logic ce12_done;
    logic [4:0] ce13_lenA;
    logic [4:0] ce13_lenB;
    logic [4:0] ce13_addrA;
    logic [4:0] ce13_addrB;
    logic ce13_mlA;
    logic ce13_mlB;
    logic [4:0] ce13_lenX;
    logic [4:0] ce13_addrX;
    logic ce13_mlX;
    logic ce13_go;
    logic ce13_clk;
    logic ce13_reset;
    logic ce13_done;
    logic [4:0] ce14_lenA;
    logic [4:0] ce14_lenB;
    logic [4:0] ce14_addrA;
    logic [4:0] ce14_addrB;
    logic ce14_mlA;
    logic ce14_mlB;
    logic [4:0] ce14_lenX;
    logic [4:0] ce14_addrX;
    logic ce14_mlX;
    logic ce14_go;
    logic ce14_clk;
    logic ce14_reset;
    logic ce14_done;
    logic [4:0] ce15_lenA;
    logic [4:0] ce15_lenB;
    logic [4:0] ce15_addrA;
    logic [4:0] ce15_addrB;
    logic ce15_mlA;
    logic ce15_mlB;
    logic [4:0] ce15_lenX;
    logic [4:0] ce15_addrX;
    logic ce15_mlX;
    logic ce15_go;
    logic ce15_clk;
    logic ce15_reset;
    logic ce15_done;
    logic [4:0] ce16_lenA;
    logic [4:0] ce16_lenB;
    logic [4:0] ce16_addrA;
    logic [4:0] ce16_addrB;
    logic ce16_mlA;
    logic ce16_mlB;
    logic [4:0] ce16_lenX;
    logic [4:0] ce16_addrX;
    logic ce16_mlX;
    logic ce16_go;
    logic ce16_clk;
    logic ce16_reset;
    logic ce16_done;
    logic [4:0] ce17_lenA;
    logic [4:0] ce17_lenB;
    logic [4:0] ce17_addrA;
    logic [4:0] ce17_addrB;
    logic ce17_mlA;
    logic ce17_mlB;
    logic [4:0] ce17_lenX;
    logic [4:0] ce17_addrX;
    logic ce17_mlX;
    logic ce17_go;
    logic ce17_clk;
    logic ce17_reset;
    logic ce17_done;
    logic [4:0] ce20_lenA;
    logic [4:0] ce20_lenB;
    logic [4:0] ce20_addrA;
    logic [4:0] ce20_addrB;
    logic ce20_mlA;
    logic ce20_mlB;
    logic [4:0] ce20_lenX;
    logic [4:0] ce20_addrX;
    logic ce20_mlX;
    logic ce20_go;
    logic ce20_clk;
    logic ce20_reset;
    logic ce20_done;
    logic [4:0] ce21_lenA;
    logic [4:0] ce21_lenB;
    logic [4:0] ce21_addrA;
    logic [4:0] ce21_addrB;
    logic ce21_mlA;
    logic ce21_mlB;
    logic [4:0] ce21_lenX;
    logic [4:0] ce21_addrX;
    logic ce21_mlX;
    logic ce21_go;
    logic ce21_clk;
    logic ce21_reset;
    logic ce21_done;
    logic [4:0] ce22_lenA;
    logic [4:0] ce22_lenB;
    logic [4:0] ce22_addrA;
    logic [4:0] ce22_addrB;
    logic ce22_mlA;
    logic ce22_mlB;
    logic [4:0] ce22_lenX;
    logic [4:0] ce22_addrX;
    logic ce22_mlX;
    logic ce22_go;
    logic ce22_clk;
    logic ce22_reset;
    logic ce22_done;
    logic [4:0] ce23_lenA;
    logic [4:0] ce23_lenB;
    logic [4:0] ce23_addrA;
    logic [4:0] ce23_addrB;
    logic ce23_mlA;
    logic ce23_mlB;
    logic [4:0] ce23_lenX;
    logic [4:0] ce23_addrX;
    logic ce23_mlX;
    logic ce23_go;
    logic ce23_clk;
    logic ce23_reset;
    logic ce23_done;
    logic [4:0] ce30_lenA;
    logic [4:0] ce30_lenB;
    logic [4:0] ce30_addrA;
    logic [4:0] ce30_addrB;
    logic ce30_mlA;
    logic ce30_mlB;
    logic [4:0] ce30_lenX;
    logic [4:0] ce30_addrX;
    logic ce30_mlX;
    logic ce30_go;
    logic ce30_clk;
    logic ce30_reset;
    logic ce30_done;
    logic [4:0] ce31_lenA;
    logic [4:0] ce31_lenB;
    logic [4:0] ce31_addrA;
    logic [4:0] ce31_addrB;
    logic ce31_mlA;
    logic ce31_mlB;
    logic [4:0] ce31_lenX;
    logic [4:0] ce31_addrX;
    logic ce31_mlX;
    logic ce31_go;
    logic ce31_clk;
    logic ce31_reset;
    logic ce31_done;
    logic [4:0] ce40_lenA;
    logic [4:0] ce40_lenB;
    logic [4:0] ce40_addrA;
    logic [4:0] ce40_addrB;
    logic ce40_mlA;
    logic ce40_mlB;
    logic [4:0] ce40_lenX;
    logic [4:0] ce40_addrX;
    logic ce40_mlX;
    logic ce40_go;
    logic ce40_clk;
    logic ce40_reset;
    logic ce40_done;
    logic comb_reg0_in;
    logic comb_reg0_write_en;
    logic comb_reg0_clk;
    logic comb_reg0_reset;
    logic comb_reg0_out;
    logic comb_reg0_done;
    logic comb_reg1_in;
    logic comb_reg1_write_en;
    logic comb_reg1_clk;
    logic comb_reg1_reset;
    logic comb_reg1_out;
    logic comb_reg1_done;
    logic comb_reg2_in;
    logic comb_reg2_write_en;
    logic comb_reg2_clk;
    logic comb_reg2_reset;
    logic comb_reg2_out;
    logic comb_reg2_done;
    logic comb_reg3_in;
    logic comb_reg3_write_en;
    logic comb_reg3_clk;
    logic comb_reg3_reset;
    logic comb_reg3_out;
    logic comb_reg3_done;
    logic comb_reg4_in;
    logic comb_reg4_write_en;
    logic comb_reg4_clk;
    logic comb_reg4_reset;
    logic comb_reg4_out;
    logic comb_reg4_done;
    logic comb_reg5_in;
    logic comb_reg5_write_en;
    logic comb_reg5_clk;
    logic comb_reg5_reset;
    logic comb_reg5_out;
    logic comb_reg5_done;
    logic comb_reg6_in;
    logic comb_reg6_write_en;
    logic comb_reg6_clk;
    logic comb_reg6_reset;
    logic comb_reg6_out;
    logic comb_reg6_done;
    logic comb_reg7_in;
    logic comb_reg7_write_en;
    logic comb_reg7_clk;
    logic comb_reg7_reset;
    logic comb_reg7_out;
    logic comb_reg7_done;
    logic comb_reg8_in;
    logic comb_reg8_write_en;
    logic comb_reg8_clk;
    logic comb_reg8_reset;
    logic comb_reg8_out;
    logic comb_reg8_done;
    logic comb_reg9_in;
    logic comb_reg9_write_en;
    logic comb_reg9_clk;
    logic comb_reg9_reset;
    logic comb_reg9_out;
    logic comb_reg9_done;
    logic comb_reg10_in;
    logic comb_reg10_write_en;
    logic comb_reg10_clk;
    logic comb_reg10_reset;
    logic comb_reg10_out;
    logic comb_reg10_done;
    logic comb_reg11_in;
    logic comb_reg11_write_en;
    logic comb_reg11_clk;
    logic comb_reg11_reset;
    logic comb_reg11_out;
    logic comb_reg11_done;
    logic comb_reg12_in;
    logic comb_reg12_write_en;
    logic comb_reg12_clk;
    logic comb_reg12_reset;
    logic comb_reg12_out;
    logic comb_reg12_done;
    logic comb_reg13_in;
    logic comb_reg13_write_en;
    logic comb_reg13_clk;
    logic comb_reg13_reset;
    logic comb_reg13_out;
    logic comb_reg13_done;
    logic comb_reg14_in;
    logic comb_reg14_write_en;
    logic comb_reg14_clk;
    logic comb_reg14_reset;
    logic comb_reg14_out;
    logic comb_reg14_done;
    logic comb_reg15_in;
    logic comb_reg15_write_en;
    logic comb_reg15_clk;
    logic comb_reg15_reset;
    logic comb_reg15_out;
    logic comb_reg15_done;
    logic comb_reg16_in;
    logic comb_reg16_write_en;
    logic comb_reg16_clk;
    logic comb_reg16_reset;
    logic comb_reg16_out;
    logic comb_reg16_done;
    logic comb_reg17_in;
    logic comb_reg17_write_en;
    logic comb_reg17_clk;
    logic comb_reg17_reset;
    logic comb_reg17_out;
    logic comb_reg17_done;
    logic comb_reg18_in;
    logic comb_reg18_write_en;
    logic comb_reg18_clk;
    logic comb_reg18_reset;
    logic comb_reg18_out;
    logic comb_reg18_done;
    logic comb_reg19_in;
    logic comb_reg19_write_en;
    logic comb_reg19_clk;
    logic comb_reg19_reset;
    logic comb_reg19_out;
    logic comb_reg19_done;
    logic comb_reg20_in;
    logic comb_reg20_write_en;
    logic comb_reg20_clk;
    logic comb_reg20_reset;
    logic comb_reg20_out;
    logic comb_reg20_done;
    logic comb_reg21_in;
    logic comb_reg21_write_en;
    logic comb_reg21_clk;
    logic comb_reg21_reset;
    logic comb_reg21_out;
    logic comb_reg21_done;
    logic comb_reg22_in;
    logic comb_reg22_write_en;
    logic comb_reg22_clk;
    logic comb_reg22_reset;
    logic comb_reg22_out;
    logic comb_reg22_done;
    logic comb_reg23_in;
    logic comb_reg23_write_en;
    logic comb_reg23_clk;
    logic comb_reg23_reset;
    logic comb_reg23_out;
    logic comb_reg23_done;
    logic comb_reg24_in;
    logic comb_reg24_write_en;
    logic comb_reg24_clk;
    logic comb_reg24_reset;
    logic comb_reg24_out;
    logic comb_reg24_done;
    logic comb_reg25_in;
    logic comb_reg25_write_en;
    logic comb_reg25_clk;
    logic comb_reg25_reset;
    logic comb_reg25_out;
    logic comb_reg25_done;
    logic comb_reg26_in;
    logic comb_reg26_write_en;
    logic comb_reg26_clk;
    logic comb_reg26_reset;
    logic comb_reg26_out;
    logic comb_reg26_done;
    logic comb_reg27_in;
    logic comb_reg27_write_en;
    logic comb_reg27_clk;
    logic comb_reg27_reset;
    logic comb_reg27_out;
    logic comb_reg27_done;
    logic comb_reg28_in;
    logic comb_reg28_write_en;
    logic comb_reg28_clk;
    logic comb_reg28_reset;
    logic comb_reg28_out;
    logic comb_reg28_done;
    logic comb_reg29_in;
    logic comb_reg29_write_en;
    logic comb_reg29_clk;
    logic comb_reg29_reset;
    logic comb_reg29_out;
    logic comb_reg29_done;
    logic comb_reg30_in;
    logic comb_reg30_write_en;
    logic comb_reg30_clk;
    logic comb_reg30_reset;
    logic comb_reg30_out;
    logic comb_reg30_done;
    logic comb_reg31_in;
    logic comb_reg31_write_en;
    logic comb_reg31_clk;
    logic comb_reg31_reset;
    logic comb_reg31_out;
    logic comb_reg31_done;
    logic [4:0] out_in;
    logic out_write_en;
    logic out_clk;
    logic out_reset;
    logic [4:0] out_out;
    logic out_done;
    logic [1:0] fsm_in;
    logic fsm_write_en;
    logic fsm_clk;
    logic fsm_reset;
    logic [1:0] fsm_out;
    logic fsm_done;
    logic pd_in;
    logic pd_write_en;
    logic pd_clk;
    logic pd_reset;
    logic pd_out;
    logic pd_done;
    logic [1:0] fsm0_in;
    logic fsm0_write_en;
    logic fsm0_clk;
    logic fsm0_reset;
    logic [1:0] fsm0_out;
    logic fsm0_done;
    logic pd0_in;
    logic pd0_write_en;
    logic pd0_clk;
    logic pd0_reset;
    logic pd0_out;
    logic pd0_done;
    logic [1:0] fsm1_in;
    logic fsm1_write_en;
    logic fsm1_clk;
    logic fsm1_reset;
    logic [1:0] fsm1_out;
    logic fsm1_done;
    logic pd1_in;
    logic pd1_write_en;
    logic pd1_clk;
    logic pd1_reset;
    logic pd1_out;
    logic pd1_done;
    logic [1:0] fsm2_in;
    logic fsm2_write_en;
    logic fsm2_clk;
    logic fsm2_reset;
    logic [1:0] fsm2_out;
    logic fsm2_done;
    logic pd2_in;
    logic pd2_write_en;
    logic pd2_clk;
    logic pd2_reset;
    logic pd2_out;
    logic pd2_done;
    logic [1:0] fsm3_in;
    logic fsm3_write_en;
    logic fsm3_clk;
    logic fsm3_reset;
    logic [1:0] fsm3_out;
    logic fsm3_done;
    logic pd3_in;
    logic pd3_write_en;
    logic pd3_clk;
    logic pd3_reset;
    logic pd3_out;
    logic pd3_done;
    logic [1:0] fsm4_in;
    logic fsm4_write_en;
    logic fsm4_clk;
    logic fsm4_reset;
    logic [1:0] fsm4_out;
    logic fsm4_done;
    logic pd4_in;
    logic pd4_write_en;
    logic pd4_clk;
    logic pd4_reset;
    logic pd4_out;
    logic pd4_done;
    logic [1:0] fsm5_in;
    logic fsm5_write_en;
    logic fsm5_clk;
    logic fsm5_reset;
    logic [1:0] fsm5_out;
    logic fsm5_done;
    logic pd5_in;
    logic pd5_write_en;
    logic pd5_clk;
    logic pd5_reset;
    logic pd5_out;
    logic pd5_done;
    logic [1:0] fsm6_in;
    logic fsm6_write_en;
    logic fsm6_clk;
    logic fsm6_reset;
    logic [1:0] fsm6_out;
    logic fsm6_done;
    logic pd6_in;
    logic pd6_write_en;
    logic pd6_clk;
    logic pd6_reset;
    logic pd6_out;
    logic pd6_done;
    logic [1:0] fsm7_in;
    logic fsm7_write_en;
    logic fsm7_clk;
    logic fsm7_reset;
    logic [1:0] fsm7_out;
    logic fsm7_done;
    logic pd7_in;
    logic pd7_write_en;
    logic pd7_clk;
    logic pd7_reset;
    logic pd7_out;
    logic pd7_done;
    logic [1:0] fsm8_in;
    logic fsm8_write_en;
    logic fsm8_clk;
    logic fsm8_reset;
    logic [1:0] fsm8_out;
    logic fsm8_done;
    logic pd8_in;
    logic pd8_write_en;
    logic pd8_clk;
    logic pd8_reset;
    logic pd8_out;
    logic pd8_done;
    logic [1:0] fsm9_in;
    logic fsm9_write_en;
    logic fsm9_clk;
    logic fsm9_reset;
    logic [1:0] fsm9_out;
    logic fsm9_done;
    logic pd9_in;
    logic pd9_write_en;
    logic pd9_clk;
    logic pd9_reset;
    logic pd9_out;
    logic pd9_done;
    logic [1:0] fsm10_in;
    logic fsm10_write_en;
    logic fsm10_clk;
    logic fsm10_reset;
    logic [1:0] fsm10_out;
    logic fsm10_done;
    logic pd10_in;
    logic pd10_write_en;
    logic pd10_clk;
    logic pd10_reset;
    logic pd10_out;
    logic pd10_done;
    logic [1:0] fsm11_in;
    logic fsm11_write_en;
    logic fsm11_clk;
    logic fsm11_reset;
    logic [1:0] fsm11_out;
    logic fsm11_done;
    logic pd11_in;
    logic pd11_write_en;
    logic pd11_clk;
    logic pd11_reset;
    logic pd11_out;
    logic pd11_done;
    logic [1:0] fsm12_in;
    logic fsm12_write_en;
    logic fsm12_clk;
    logic fsm12_reset;
    logic [1:0] fsm12_out;
    logic fsm12_done;
    logic pd12_in;
    logic pd12_write_en;
    logic pd12_clk;
    logic pd12_reset;
    logic pd12_out;
    logic pd12_done;
    logic [1:0] fsm13_in;
    logic fsm13_write_en;
    logic fsm13_clk;
    logic fsm13_reset;
    logic [1:0] fsm13_out;
    logic fsm13_done;
    logic pd13_in;
    logic pd13_write_en;
    logic pd13_clk;
    logic pd13_reset;
    logic pd13_out;
    logic pd13_done;
    logic [1:0] fsm14_in;
    logic fsm14_write_en;
    logic fsm14_clk;
    logic fsm14_reset;
    logic [1:0] fsm14_out;
    logic fsm14_done;
    logic pd14_in;
    logic pd14_write_en;
    logic pd14_clk;
    logic pd14_reset;
    logic pd14_out;
    logic pd14_done;
    logic [1:0] fsm15_in;
    logic fsm15_write_en;
    logic fsm15_clk;
    logic fsm15_reset;
    logic [1:0] fsm15_out;
    logic fsm15_done;
    logic pd15_in;
    logic pd15_write_en;
    logic pd15_clk;
    logic pd15_reset;
    logic pd15_out;
    logic pd15_done;
    logic [1:0] fsm16_in;
    logic fsm16_write_en;
    logic fsm16_clk;
    logic fsm16_reset;
    logic [1:0] fsm16_out;
    logic fsm16_done;
    logic pd16_in;
    logic pd16_write_en;
    logic pd16_clk;
    logic pd16_reset;
    logic pd16_out;
    logic pd16_done;
    logic [1:0] fsm17_in;
    logic fsm17_write_en;
    logic fsm17_clk;
    logic fsm17_reset;
    logic [1:0] fsm17_out;
    logic fsm17_done;
    logic pd17_in;
    logic pd17_write_en;
    logic pd17_clk;
    logic pd17_reset;
    logic pd17_out;
    logic pd17_done;
    logic [1:0] fsm18_in;
    logic fsm18_write_en;
    logic fsm18_clk;
    logic fsm18_reset;
    logic [1:0] fsm18_out;
    logic fsm18_done;
    logic pd18_in;
    logic pd18_write_en;
    logic pd18_clk;
    logic pd18_reset;
    logic pd18_out;
    logic pd18_done;
    logic [1:0] fsm19_in;
    logic fsm19_write_en;
    logic fsm19_clk;
    logic fsm19_reset;
    logic [1:0] fsm19_out;
    logic fsm19_done;
    logic pd19_in;
    logic pd19_write_en;
    logic pd19_clk;
    logic pd19_reset;
    logic pd19_out;
    logic pd19_done;
    logic [1:0] fsm20_in;
    logic fsm20_write_en;
    logic fsm20_clk;
    logic fsm20_reset;
    logic [1:0] fsm20_out;
    logic fsm20_done;
    logic pd20_in;
    logic pd20_write_en;
    logic pd20_clk;
    logic pd20_reset;
    logic pd20_out;
    logic pd20_done;
    logic [1:0] fsm21_in;
    logic fsm21_write_en;
    logic fsm21_clk;
    logic fsm21_reset;
    logic [1:0] fsm21_out;
    logic fsm21_done;
    logic pd21_in;
    logic pd21_write_en;
    logic pd21_clk;
    logic pd21_reset;
    logic pd21_out;
    logic pd21_done;
    logic [1:0] fsm22_in;
    logic fsm22_write_en;
    logic fsm22_clk;
    logic fsm22_reset;
    logic [1:0] fsm22_out;
    logic fsm22_done;
    logic pd22_in;
    logic pd22_write_en;
    logic pd22_clk;
    logic pd22_reset;
    logic pd22_out;
    logic pd22_done;
    logic [1:0] fsm23_in;
    logic fsm23_write_en;
    logic fsm23_clk;
    logic fsm23_reset;
    logic [1:0] fsm23_out;
    logic fsm23_done;
    logic pd23_in;
    logic pd23_write_en;
    logic pd23_clk;
    logic pd23_reset;
    logic pd23_out;
    logic pd23_done;
    logic [1:0] fsm24_in;
    logic fsm24_write_en;
    logic fsm24_clk;
    logic fsm24_reset;
    logic [1:0] fsm24_out;
    logic fsm24_done;
    logic pd24_in;
    logic pd24_write_en;
    logic pd24_clk;
    logic pd24_reset;
    logic pd24_out;
    logic pd24_done;
    logic [1:0] fsm25_in;
    logic fsm25_write_en;
    logic fsm25_clk;
    logic fsm25_reset;
    logic [1:0] fsm25_out;
    logic fsm25_done;
    logic pd25_in;
    logic pd25_write_en;
    logic pd25_clk;
    logic pd25_reset;
    logic pd25_out;
    logic pd25_done;
    logic [1:0] fsm26_in;
    logic fsm26_write_en;
    logic fsm26_clk;
    logic fsm26_reset;
    logic [1:0] fsm26_out;
    logic fsm26_done;
    logic pd26_in;
    logic pd26_write_en;
    logic pd26_clk;
    logic pd26_reset;
    logic pd26_out;
    logic pd26_done;
    logic [1:0] fsm27_in;
    logic fsm27_write_en;
    logic fsm27_clk;
    logic fsm27_reset;
    logic [1:0] fsm27_out;
    logic fsm27_done;
    logic pd27_in;
    logic pd27_write_en;
    logic pd27_clk;
    logic pd27_reset;
    logic pd27_out;
    logic pd27_done;
    logic [1:0] fsm28_in;
    logic fsm28_write_en;
    logic fsm28_clk;
    logic fsm28_reset;
    logic [1:0] fsm28_out;
    logic fsm28_done;
    logic pd28_in;
    logic pd28_write_en;
    logic pd28_clk;
    logic pd28_reset;
    logic pd28_out;
    logic pd28_done;
    logic [1:0] fsm29_in;
    logic fsm29_write_en;
    logic fsm29_clk;
    logic fsm29_reset;
    logic [1:0] fsm29_out;
    logic fsm29_done;
    logic pd29_in;
    logic pd29_write_en;
    logic pd29_clk;
    logic pd29_reset;
    logic pd29_out;
    logic pd29_done;
    logic [1:0] fsm30_in;
    logic fsm30_write_en;
    logic fsm30_clk;
    logic fsm30_reset;
    logic [1:0] fsm30_out;
    logic fsm30_done;
    logic pd30_in;
    logic pd30_write_en;
    logic pd30_clk;
    logic pd30_reset;
    logic pd30_out;
    logic pd30_done;
    logic pd31_in;
    logic pd31_write_en;
    logic pd31_clk;
    logic pd31_reset;
    logic pd31_out;
    logic pd31_done;
    logic pd32_in;
    logic pd32_write_en;
    logic pd32_clk;
    logic pd32_reset;
    logic pd32_out;
    logic pd32_done;
    logic pd33_in;
    logic pd33_write_en;
    logic pd33_clk;
    logic pd33_reset;
    logic pd33_out;
    logic pd33_done;
    logic pd34_in;
    logic pd34_write_en;
    logic pd34_clk;
    logic pd34_reset;
    logic pd34_out;
    logic pd34_done;
    logic pd35_in;
    logic pd35_write_en;
    logic pd35_clk;
    logic pd35_reset;
    logic pd35_out;
    logic pd35_done;
    logic pd36_in;
    logic pd36_write_en;
    logic pd36_clk;
    logic pd36_reset;
    logic pd36_out;
    logic pd36_done;
    logic pd37_in;
    logic pd37_write_en;
    logic pd37_clk;
    logic pd37_reset;
    logic pd37_out;
    logic pd37_done;
    logic pd38_in;
    logic pd38_write_en;
    logic pd38_clk;
    logic pd38_reset;
    logic pd38_out;
    logic pd38_done;
    logic pd39_in;
    logic pd39_write_en;
    logic pd39_clk;
    logic pd39_reset;
    logic pd39_out;
    logic pd39_done;
    logic pd40_in;
    logic pd40_write_en;
    logic pd40_clk;
    logic pd40_reset;
    logic pd40_out;
    logic pd40_done;
    logic pd41_in;
    logic pd41_write_en;
    logic pd41_clk;
    logic pd41_reset;
    logic pd41_out;
    logic pd41_done;
    logic pd42_in;
    logic pd42_write_en;
    logic pd42_clk;
    logic pd42_reset;
    logic pd42_out;
    logic pd42_done;
    logic pd43_in;
    logic pd43_write_en;
    logic pd43_clk;
    logic pd43_reset;
    logic pd43_out;
    logic pd43_done;
    logic pd44_in;
    logic pd44_write_en;
    logic pd44_clk;
    logic pd44_reset;
    logic pd44_out;
    logic pd44_done;
    logic pd45_in;
    logic pd45_write_en;
    logic pd45_clk;
    logic pd45_reset;
    logic pd45_out;
    logic pd45_done;
    logic pd46_in;
    logic pd46_write_en;
    logic pd46_clk;
    logic pd46_reset;
    logic pd46_out;
    logic pd46_done;
    logic pd47_in;
    logic pd47_write_en;
    logic pd47_clk;
    logic pd47_reset;
    logic pd47_out;
    logic pd47_done;
    logic pd48_in;
    logic pd48_write_en;
    logic pd48_clk;
    logic pd48_reset;
    logic pd48_out;
    logic pd48_done;
    logic pd49_in;
    logic pd49_write_en;
    logic pd49_clk;
    logic pd49_reset;
    logic pd49_out;
    logic pd49_done;
    logic pd50_in;
    logic pd50_write_en;
    logic pd50_clk;
    logic pd50_reset;
    logic pd50_out;
    logic pd50_done;
    logic pd51_in;
    logic pd51_write_en;
    logic pd51_clk;
    logic pd51_reset;
    logic pd51_out;
    logic pd51_done;
    logic pd52_in;
    logic pd52_write_en;
    logic pd52_clk;
    logic pd52_reset;
    logic pd52_out;
    logic pd52_done;
    logic pd53_in;
    logic pd53_write_en;
    logic pd53_clk;
    logic pd53_reset;
    logic pd53_out;
    logic pd53_done;
    logic pd54_in;
    logic pd54_write_en;
    logic pd54_clk;
    logic pd54_reset;
    logic pd54_out;
    logic pd54_done;
    logic pd55_in;
    logic pd55_write_en;
    logic pd55_clk;
    logic pd55_reset;
    logic pd55_out;
    logic pd55_done;
    logic pd56_in;
    logic pd56_write_en;
    logic pd56_clk;
    logic pd56_reset;
    logic pd56_out;
    logic pd56_done;
    logic pd57_in;
    logic pd57_write_en;
    logic pd57_clk;
    logic pd57_reset;
    logic pd57_out;
    logic pd57_done;
    logic pd58_in;
    logic pd58_write_en;
    logic pd58_clk;
    logic pd58_reset;
    logic pd58_out;
    logic pd58_done;
    logic pd59_in;
    logic pd59_write_en;
    logic pd59_clk;
    logic pd59_reset;
    logic pd59_out;
    logic pd59_done;
    logic pd60_in;
    logic pd60_write_en;
    logic pd60_clk;
    logic pd60_reset;
    logic pd60_out;
    logic pd60_done;
    logic pd61_in;
    logic pd61_write_en;
    logic pd61_clk;
    logic pd61_reset;
    logic pd61_out;
    logic pd61_done;
    logic pd62_in;
    logic pd62_write_en;
    logic pd62_clk;
    logic pd62_reset;
    logic pd62_out;
    logic pd62_done;
    logic pd63_in;
    logic pd63_write_en;
    logic pd63_clk;
    logic pd63_reset;
    logic pd63_out;
    logic pd63_done;
    logic pd64_in;
    logic pd64_write_en;
    logic pd64_clk;
    logic pd64_reset;
    logic pd64_out;
    logic pd64_done;
    logic pd65_in;
    logic pd65_write_en;
    logic pd65_clk;
    logic pd65_reset;
    logic pd65_out;
    logic pd65_done;
    logic pd66_in;
    logic pd66_write_en;
    logic pd66_clk;
    logic pd66_reset;
    logic pd66_out;
    logic pd66_done;
    logic pd67_in;
    logic pd67_write_en;
    logic pd67_clk;
    logic pd67_reset;
    logic pd67_out;
    logic pd67_done;
    logic pd68_in;
    logic pd68_write_en;
    logic pd68_clk;
    logic pd68_reset;
    logic pd68_out;
    logic pd68_done;
    logic pd69_in;
    logic pd69_write_en;
    logic pd69_clk;
    logic pd69_reset;
    logic pd69_out;
    logic pd69_done;
    logic pd70_in;
    logic pd70_write_en;
    logic pd70_clk;
    logic pd70_reset;
    logic pd70_out;
    logic pd70_done;
    logic pd71_in;
    logic pd71_write_en;
    logic pd71_clk;
    logic pd71_reset;
    logic pd71_out;
    logic pd71_done;
    logic pd72_in;
    logic pd72_write_en;
    logic pd72_clk;
    logic pd72_reset;
    logic pd72_out;
    logic pd72_done;
    logic pd73_in;
    logic pd73_write_en;
    logic pd73_clk;
    logic pd73_reset;
    logic pd73_out;
    logic pd73_done;
    logic pd74_in;
    logic pd74_write_en;
    logic pd74_clk;
    logic pd74_reset;
    logic pd74_out;
    logic pd74_done;
    logic pd75_in;
    logic pd75_write_en;
    logic pd75_clk;
    logic pd75_reset;
    logic pd75_out;
    logic pd75_done;
    logic pd76_in;
    logic pd76_write_en;
    logic pd76_clk;
    logic pd76_reset;
    logic pd76_out;
    logic pd76_done;
    logic pd77_in;
    logic pd77_write_en;
    logic pd77_clk;
    logic pd77_reset;
    logic pd77_out;
    logic pd77_done;
    logic pd78_in;
    logic pd78_write_en;
    logic pd78_clk;
    logic pd78_reset;
    logic pd78_out;
    logic pd78_done;
    logic pd79_in;
    logic pd79_write_en;
    logic pd79_clk;
    logic pd79_reset;
    logic pd79_out;
    logic pd79_done;
    logic pd80_in;
    logic pd80_write_en;
    logic pd80_clk;
    logic pd80_reset;
    logic pd80_out;
    logic pd80_done;
    logic pd81_in;
    logic pd81_write_en;
    logic pd81_clk;
    logic pd81_reset;
    logic pd81_out;
    logic pd81_done;
    logic pd82_in;
    logic pd82_write_en;
    logic pd82_clk;
    logic pd82_reset;
    logic pd82_out;
    logic pd82_done;
    logic pd83_in;
    logic pd83_write_en;
    logic pd83_clk;
    logic pd83_reset;
    logic pd83_out;
    logic pd83_done;
    logic pd84_in;
    logic pd84_write_en;
    logic pd84_clk;
    logic pd84_reset;
    logic pd84_out;
    logic pd84_done;
    logic pd85_in;
    logic pd85_write_en;
    logic pd85_clk;
    logic pd85_reset;
    logic pd85_out;
    logic pd85_done;
    logic pd86_in;
    logic pd86_write_en;
    logic pd86_clk;
    logic pd86_reset;
    logic pd86_out;
    logic pd86_done;
    logic pd87_in;
    logic pd87_write_en;
    logic pd87_clk;
    logic pd87_reset;
    logic pd87_out;
    logic pd87_done;
    logic pd88_in;
    logic pd88_write_en;
    logic pd88_clk;
    logic pd88_reset;
    logic pd88_out;
    logic pd88_done;
    logic pd89_in;
    logic pd89_write_en;
    logic pd89_clk;
    logic pd89_reset;
    logic pd89_out;
    logic pd89_done;
    logic pd90_in;
    logic pd90_write_en;
    logic pd90_clk;
    logic pd90_reset;
    logic pd90_out;
    logic pd90_done;
    logic pd91_in;
    logic pd91_write_en;
    logic pd91_clk;
    logic pd91_reset;
    logic pd91_out;
    logic pd91_done;
    logic pd92_in;
    logic pd92_write_en;
    logic pd92_clk;
    logic pd92_reset;
    logic pd92_out;
    logic pd92_done;
    logic [2:0] fsm31_in;
    logic fsm31_write_en;
    logic fsm31_clk;
    logic fsm31_reset;
    logic [2:0] fsm31_out;
    logic fsm31_done;
    logic pd93_in;
    logic pd93_write_en;
    logic pd93_clk;
    logic pd93_reset;
    logic pd93_out;
    logic pd93_done;
    logic [3:0] fsm32_in;
    logic fsm32_write_en;
    logic fsm32_clk;
    logic fsm32_reset;
    logic [3:0] fsm32_out;
    logic fsm32_done;
    logic pd94_in;
    logic pd94_write_en;
    logic pd94_clk;
    logic pd94_reset;
    logic pd94_out;
    logic pd94_done;
    logic fsm33_in;
    logic fsm33_write_en;
    logic fsm33_clk;
    logic fsm33_reset;
    logic fsm33_out;
    logic fsm33_done;
    logic write_zero_go_in;
    logic write_zero_go_out;
    logic write_zero_done_in;
    logic write_zero_done_out;
    logic write0_go_in;
    logic write0_go_out;
    logic write0_done_in;
    logic write0_done_out;
    logic write1_go_in;
    logic write1_go_out;
    logic write1_done_in;
    logic write1_done_out;
    logic write2_go_in;
    logic write2_go_out;
    logic write2_done_in;
    logic write2_done_out;
    logic write3_go_in;
    logic write3_go_out;
    logic write3_done_in;
    logic write3_done_out;
    logic write4_go_in;
    logic write4_go_out;
    logic write4_done_in;
    logic write4_done_out;
    logic write5_go_in;
    logic write5_go_out;
    logic write5_done_in;
    logic write5_done_out;
    logic write6_go_in;
    logic write6_go_out;
    logic write6_done_in;
    logic write6_done_out;
    logic write7_go_in;
    logic write7_go_out;
    logic write7_done_in;
    logic write7_done_out;
    logic write8_go_in;
    logic write8_go_out;
    logic write8_done_in;
    logic write8_done_out;
    logic write9_go_in;
    logic write9_go_out;
    logic write9_done_in;
    logic write9_done_out;
    logic write10_go_in;
    logic write10_go_out;
    logic write10_done_in;
    logic write10_done_out;
    logic write11_go_in;
    logic write11_go_out;
    logic write11_done_in;
    logic write11_done_out;
    logic write12_go_in;
    logic write12_go_out;
    logic write12_done_in;
    logic write12_done_out;
    logic write13_go_in;
    logic write13_go_out;
    logic write13_done_in;
    logic write13_done_out;
    logic write14_go_in;
    logic write14_go_out;
    logic write14_done_in;
    logic write14_done_out;
    logic write15_go_in;
    logic write15_go_out;
    logic write15_done_in;
    logic write15_done_out;
    logic write16_go_in;
    logic write16_go_out;
    logic write16_done_in;
    logic write16_done_out;
    logic write17_go_in;
    logic write17_go_out;
    logic write17_done_in;
    logic write17_done_out;
    logic write18_go_in;
    logic write18_go_out;
    logic write18_done_in;
    logic write18_done_out;
    logic write19_go_in;
    logic write19_go_out;
    logic write19_done_in;
    logic write19_done_out;
    logic write20_go_in;
    logic write20_go_out;
    logic write20_done_in;
    logic write20_done_out;
    logic write21_go_in;
    logic write21_go_out;
    logic write21_done_in;
    logic write21_done_out;
    logic write22_go_in;
    logic write22_go_out;
    logic write22_done_in;
    logic write22_done_out;
    logic write23_go_in;
    logic write23_go_out;
    logic write23_done_in;
    logic write23_done_out;
    logic write24_go_in;
    logic write24_go_out;
    logic write24_done_in;
    logic write24_done_out;
    logic write25_go_in;
    logic write25_go_out;
    logic write25_done_in;
    logic write25_done_out;
    logic write26_go_in;
    logic write26_go_out;
    logic write26_done_in;
    logic write26_done_out;
    logic write27_go_in;
    logic write27_go_out;
    logic write27_done_in;
    logic write27_done_out;
    logic write28_go_in;
    logic write28_go_out;
    logic write28_done_in;
    logic write28_done_out;
    logic write29_go_in;
    logic write29_go_out;
    logic write29_done_in;
    logic write29_done_out;
    logic write30_go_in;
    logic write30_go_out;
    logic write30_done_in;
    logic write30_done_out;
    logic write31_go_in;
    logic write31_go_out;
    logic write31_done_in;
    logic write31_done_out;
    logic find_write_index_go_in;
    logic find_write_index_go_out;
    logic find_write_index_done_in;
    logic find_write_index_done_out;
    logic default_to_zero_length_index_go_in;
    logic default_to_zero_length_index_go_out;
    logic default_to_zero_length_index_done_in;
    logic default_to_zero_length_index_done_out;
    logic save_index_go_in;
    logic save_index_go_out;
    logic save_index_done_in;
    logic save_index_done_out;
    logic is_length_zero0_go_in;
    logic is_length_zero0_go_out;
    logic is_length_zero0_done_in;
    logic is_length_zero0_done_out;
    logic invoke_go_in;
    logic invoke_go_out;
    logic invoke_done_in;
    logic invoke_done_out;
    logic invoke0_go_in;
    logic invoke0_go_out;
    logic invoke0_done_in;
    logic invoke0_done_out;
    logic invoke1_go_in;
    logic invoke1_go_out;
    logic invoke1_done_in;
    logic invoke1_done_out;
    logic invoke2_go_in;
    logic invoke2_go_out;
    logic invoke2_done_in;
    logic invoke2_done_out;
    logic invoke3_go_in;
    logic invoke3_go_out;
    logic invoke3_done_in;
    logic invoke3_done_out;
    logic invoke4_go_in;
    logic invoke4_go_out;
    logic invoke4_done_in;
    logic invoke4_done_out;
    logic invoke5_go_in;
    logic invoke5_go_out;
    logic invoke5_done_in;
    logic invoke5_done_out;
    logic invoke6_go_in;
    logic invoke6_go_out;
    logic invoke6_done_in;
    logic invoke6_done_out;
    logic invoke7_go_in;
    logic invoke7_go_out;
    logic invoke7_done_in;
    logic invoke7_done_out;
    logic invoke8_go_in;
    logic invoke8_go_out;
    logic invoke8_done_in;
    logic invoke8_done_out;
    logic invoke9_go_in;
    logic invoke9_go_out;
    logic invoke9_done_in;
    logic invoke9_done_out;
    logic invoke10_go_in;
    logic invoke10_go_out;
    logic invoke10_done_in;
    logic invoke10_done_out;
    logic invoke11_go_in;
    logic invoke11_go_out;
    logic invoke11_done_in;
    logic invoke11_done_out;
    logic invoke12_go_in;
    logic invoke12_go_out;
    logic invoke12_done_in;
    logic invoke12_done_out;
    logic invoke13_go_in;
    logic invoke13_go_out;
    logic invoke13_done_in;
    logic invoke13_done_out;
    logic invoke14_go_in;
    logic invoke14_go_out;
    logic invoke14_done_in;
    logic invoke14_done_out;
    logic invoke15_go_in;
    logic invoke15_go_out;
    logic invoke15_done_in;
    logic invoke15_done_out;
    logic invoke16_go_in;
    logic invoke16_go_out;
    logic invoke16_done_in;
    logic invoke16_done_out;
    logic invoke17_go_in;
    logic invoke17_go_out;
    logic invoke17_done_in;
    logic invoke17_done_out;
    logic invoke18_go_in;
    logic invoke18_go_out;
    logic invoke18_done_in;
    logic invoke18_done_out;
    logic invoke19_go_in;
    logic invoke19_go_out;
    logic invoke19_done_in;
    logic invoke19_done_out;
    logic invoke20_go_in;
    logic invoke20_go_out;
    logic invoke20_done_in;
    logic invoke20_done_out;
    logic invoke21_go_in;
    logic invoke21_go_out;
    logic invoke21_done_in;
    logic invoke21_done_out;
    logic invoke22_go_in;
    logic invoke22_go_out;
    logic invoke22_done_in;
    logic invoke22_done_out;
    logic invoke23_go_in;
    logic invoke23_go_out;
    logic invoke23_done_in;
    logic invoke23_done_out;
    logic invoke24_go_in;
    logic invoke24_go_out;
    logic invoke24_done_in;
    logic invoke24_done_out;
    logic invoke25_go_in;
    logic invoke25_go_out;
    logic invoke25_done_in;
    logic invoke25_done_out;
    logic invoke26_go_in;
    logic invoke26_go_out;
    logic invoke26_done_in;
    logic invoke26_done_out;
    logic invoke27_go_in;
    logic invoke27_go_out;
    logic invoke27_done_in;
    logic invoke27_done_out;
    logic invoke28_go_in;
    logic invoke28_go_out;
    logic invoke28_done_in;
    logic invoke28_done_out;
    logic invoke29_go_in;
    logic invoke29_go_out;
    logic invoke29_done_in;
    logic invoke29_done_out;
    logic invoke30_go_in;
    logic invoke30_go_out;
    logic invoke30_done_in;
    logic invoke30_done_out;
    logic invoke31_go_in;
    logic invoke31_go_out;
    logic invoke31_done_in;
    logic invoke31_done_out;
    logic invoke32_go_in;
    logic invoke32_go_out;
    logic invoke32_done_in;
    logic invoke32_done_out;
    logic invoke33_go_in;
    logic invoke33_go_out;
    logic invoke33_done_in;
    logic invoke33_done_out;
    logic invoke34_go_in;
    logic invoke34_go_out;
    logic invoke34_done_in;
    logic invoke34_done_out;
    logic invoke35_go_in;
    logic invoke35_go_out;
    logic invoke35_done_in;
    logic invoke35_done_out;
    logic invoke36_go_in;
    logic invoke36_go_out;
    logic invoke36_done_in;
    logic invoke36_done_out;
    logic invoke37_go_in;
    logic invoke37_go_out;
    logic invoke37_done_in;
    logic invoke37_done_out;
    logic invoke38_go_in;
    logic invoke38_go_out;
    logic invoke38_done_in;
    logic invoke38_done_out;
    logic invoke39_go_in;
    logic invoke39_go_out;
    logic invoke39_done_in;
    logic invoke39_done_out;
    logic invoke40_go_in;
    logic invoke40_go_out;
    logic invoke40_done_in;
    logic invoke40_done_out;
    logic invoke41_go_in;
    logic invoke41_go_out;
    logic invoke41_done_in;
    logic invoke41_done_out;
    logic invoke42_go_in;
    logic invoke42_go_out;
    logic invoke42_done_in;
    logic invoke42_done_out;
    logic invoke43_go_in;
    logic invoke43_go_out;
    logic invoke43_done_in;
    logic invoke43_done_out;
    logic invoke44_go_in;
    logic invoke44_go_out;
    logic invoke44_done_in;
    logic invoke44_done_out;
    logic invoke45_go_in;
    logic invoke45_go_out;
    logic invoke45_done_in;
    logic invoke45_done_out;
    logic invoke46_go_in;
    logic invoke46_go_out;
    logic invoke46_done_in;
    logic invoke46_done_out;
    logic invoke47_go_in;
    logic invoke47_go_out;
    logic invoke47_done_in;
    logic invoke47_done_out;
    logic invoke48_go_in;
    logic invoke48_go_out;
    logic invoke48_done_in;
    logic invoke48_done_out;
    logic invoke49_go_in;
    logic invoke49_go_out;
    logic invoke49_done_in;
    logic invoke49_done_out;
    logic invoke50_go_in;
    logic invoke50_go_out;
    logic invoke50_done_in;
    logic invoke50_done_out;
    logic invoke51_go_in;
    logic invoke51_go_out;
    logic invoke51_done_in;
    logic invoke51_done_out;
    logic invoke52_go_in;
    logic invoke52_go_out;
    logic invoke52_done_in;
    logic invoke52_done_out;
    logic invoke53_go_in;
    logic invoke53_go_out;
    logic invoke53_done_in;
    logic invoke53_done_out;
    logic invoke54_go_in;
    logic invoke54_go_out;
    logic invoke54_done_in;
    logic invoke54_done_out;
    logic invoke55_go_in;
    logic invoke55_go_out;
    logic invoke55_done_in;
    logic invoke55_done_out;
    logic invoke56_go_in;
    logic invoke56_go_out;
    logic invoke56_done_in;
    logic invoke56_done_out;
    logic invoke57_go_in;
    logic invoke57_go_out;
    logic invoke57_done_in;
    logic invoke57_done_out;
    logic invoke58_go_in;
    logic invoke58_go_out;
    logic invoke58_done_in;
    logic invoke58_done_out;
    logic invoke59_go_in;
    logic invoke59_go_out;
    logic invoke59_done_in;
    logic invoke59_done_out;
    logic invoke60_go_in;
    logic invoke60_go_out;
    logic invoke60_done_in;
    logic invoke60_done_out;
    logic invoke61_go_in;
    logic invoke61_go_out;
    logic invoke61_done_in;
    logic invoke61_done_out;
    logic par_go_in;
    logic par_go_out;
    logic par_done_in;
    logic par_done_out;
    logic tdcc_go_in;
    logic tdcc_go_out;
    logic tdcc_done_in;
    logic tdcc_done_out;
    logic tdcc0_go_in;
    logic tdcc0_go_out;
    logic tdcc0_done_in;
    logic tdcc0_done_out;
    logic tdcc1_go_in;
    logic tdcc1_go_out;
    logic tdcc1_done_in;
    logic tdcc1_done_out;
    logic tdcc2_go_in;
    logic tdcc2_go_out;
    logic tdcc2_done_in;
    logic tdcc2_done_out;
    logic tdcc3_go_in;
    logic tdcc3_go_out;
    logic tdcc3_done_in;
    logic tdcc3_done_out;
    logic tdcc4_go_in;
    logic tdcc4_go_out;
    logic tdcc4_done_in;
    logic tdcc4_done_out;
    logic tdcc5_go_in;
    logic tdcc5_go_out;
    logic tdcc5_done_in;
    logic tdcc5_done_out;
    logic tdcc6_go_in;
    logic tdcc6_go_out;
    logic tdcc6_done_in;
    logic tdcc6_done_out;
    logic tdcc7_go_in;
    logic tdcc7_go_out;
    logic tdcc7_done_in;
    logic tdcc7_done_out;
    logic tdcc8_go_in;
    logic tdcc8_go_out;
    logic tdcc8_done_in;
    logic tdcc8_done_out;
    logic tdcc9_go_in;
    logic tdcc9_go_out;
    logic tdcc9_done_in;
    logic tdcc9_done_out;
    logic tdcc10_go_in;
    logic tdcc10_go_out;
    logic tdcc10_done_in;
    logic tdcc10_done_out;
    logic tdcc11_go_in;
    logic tdcc11_go_out;
    logic tdcc11_done_in;
    logic tdcc11_done_out;
    logic tdcc12_go_in;
    logic tdcc12_go_out;
    logic tdcc12_done_in;
    logic tdcc12_done_out;
    logic tdcc13_go_in;
    logic tdcc13_go_out;
    logic tdcc13_done_in;
    logic tdcc13_done_out;
    logic tdcc14_go_in;
    logic tdcc14_go_out;
    logic tdcc14_done_in;
    logic tdcc14_done_out;
    logic tdcc15_go_in;
    logic tdcc15_go_out;
    logic tdcc15_done_in;
    logic tdcc15_done_out;
    logic tdcc16_go_in;
    logic tdcc16_go_out;
    logic tdcc16_done_in;
    logic tdcc16_done_out;
    logic tdcc17_go_in;
    logic tdcc17_go_out;
    logic tdcc17_done_in;
    logic tdcc17_done_out;
    logic tdcc18_go_in;
    logic tdcc18_go_out;
    logic tdcc18_done_in;
    logic tdcc18_done_out;
    logic tdcc19_go_in;
    logic tdcc19_go_out;
    logic tdcc19_done_in;
    logic tdcc19_done_out;
    logic tdcc20_go_in;
    logic tdcc20_go_out;
    logic tdcc20_done_in;
    logic tdcc20_done_out;
    logic tdcc21_go_in;
    logic tdcc21_go_out;
    logic tdcc21_done_in;
    logic tdcc21_done_out;
    logic tdcc22_go_in;
    logic tdcc22_go_out;
    logic tdcc22_done_in;
    logic tdcc22_done_out;
    logic tdcc23_go_in;
    logic tdcc23_go_out;
    logic tdcc23_done_in;
    logic tdcc23_done_out;
    logic tdcc24_go_in;
    logic tdcc24_go_out;
    logic tdcc24_done_in;
    logic tdcc24_done_out;
    logic tdcc25_go_in;
    logic tdcc25_go_out;
    logic tdcc25_done_in;
    logic tdcc25_done_out;
    logic tdcc26_go_in;
    logic tdcc26_go_out;
    logic tdcc26_done_in;
    logic tdcc26_done_out;
    logic tdcc27_go_in;
    logic tdcc27_go_out;
    logic tdcc27_done_in;
    logic tdcc27_done_out;
    logic tdcc28_go_in;
    logic tdcc28_go_out;
    logic tdcc28_done_in;
    logic tdcc28_done_out;
    logic tdcc29_go_in;
    logic tdcc29_go_out;
    logic tdcc29_done_in;
    logic tdcc29_done_out;
    logic tdcc30_go_in;
    logic tdcc30_go_out;
    logic tdcc30_done_in;
    logic tdcc30_done_out;
    logic par0_go_in;
    logic par0_go_out;
    logic par0_done_in;
    logic par0_done_out;
    logic par1_go_in;
    logic par1_go_out;
    logic par1_done_in;
    logic par1_done_out;
    logic par2_go_in;
    logic par2_go_out;
    logic par2_done_in;
    logic par2_done_out;
    logic par3_go_in;
    logic par3_go_out;
    logic par3_done_in;
    logic par3_done_out;
    logic par4_go_in;
    logic par4_go_out;
    logic par4_done_in;
    logic par4_done_out;
    logic par5_go_in;
    logic par5_go_out;
    logic par5_done_in;
    logic par5_done_out;
    logic tdcc31_go_in;
    logic tdcc31_go_out;
    logic tdcc31_done_in;
    logic tdcc31_done_out;
    logic tdcc32_go_in;
    logic tdcc32_go_out;
    logic tdcc32_done_in;
    logic tdcc32_done_out;
    logic tdcc33_go_in;
    logic tdcc33_go_out;
    logic tdcc33_done_in;
    logic tdcc33_done_out;
    initial begin
        p0_in = 32'd0;
        p0_write_en = 1'd0;
        p0_clk = 1'd0;
        p0_reset = 1'd0;
        p1_in = 32'd0;
        p1_write_en = 1'd0;
        p1_clk = 1'd0;
        p1_reset = 1'd0;
        p2_in = 32'd0;
        p2_write_en = 1'd0;
        p2_clk = 1'd0;
        p2_reset = 1'd0;
        p3_in = 32'd0;
        p3_write_en = 1'd0;
        p3_clk = 1'd0;
        p3_reset = 1'd0;
        p4_in = 32'd0;
        p4_write_en = 1'd0;
        p4_clk = 1'd0;
        p4_reset = 1'd0;
        p5_in = 32'd0;
        p5_write_en = 1'd0;
        p5_clk = 1'd0;
        p5_reset = 1'd0;
        p6_in = 32'd0;
        p6_write_en = 1'd0;
        p6_clk = 1'd0;
        p6_reset = 1'd0;
        p7_in = 32'd0;
        p7_write_en = 1'd0;
        p7_clk = 1'd0;
        p7_reset = 1'd0;
        p8_in = 32'd0;
        p8_write_en = 1'd0;
        p8_clk = 1'd0;
        p8_reset = 1'd0;
        p9_in = 32'd0;
        p9_write_en = 1'd0;
        p9_clk = 1'd0;
        p9_reset = 1'd0;
        p10_in = 32'd0;
        p10_write_en = 1'd0;
        p10_clk = 1'd0;
        p10_reset = 1'd0;
        p11_in = 32'd0;
        p11_write_en = 1'd0;
        p11_clk = 1'd0;
        p11_reset = 1'd0;
        p12_in = 32'd0;
        p12_write_en = 1'd0;
        p12_clk = 1'd0;
        p12_reset = 1'd0;
        p13_in = 32'd0;
        p13_write_en = 1'd0;
        p13_clk = 1'd0;
        p13_reset = 1'd0;
        p14_in = 32'd0;
        p14_write_en = 1'd0;
        p14_clk = 1'd0;
        p14_reset = 1'd0;
        p15_in = 32'd0;
        p15_write_en = 1'd0;
        p15_clk = 1'd0;
        p15_reset = 1'd0;
        p16_in = 32'd0;
        p16_write_en = 1'd0;
        p16_clk = 1'd0;
        p16_reset = 1'd0;
        p17_in = 32'd0;
        p17_write_en = 1'd0;
        p17_clk = 1'd0;
        p17_reset = 1'd0;
        p18_in = 32'd0;
        p18_write_en = 1'd0;
        p18_clk = 1'd0;
        p18_reset = 1'd0;
        p19_in = 32'd0;
        p19_write_en = 1'd0;
        p19_clk = 1'd0;
        p19_reset = 1'd0;
        p20_in = 32'd0;
        p20_write_en = 1'd0;
        p20_clk = 1'd0;
        p20_reset = 1'd0;
        p21_in = 32'd0;
        p21_write_en = 1'd0;
        p21_clk = 1'd0;
        p21_reset = 1'd0;
        p22_in = 32'd0;
        p22_write_en = 1'd0;
        p22_clk = 1'd0;
        p22_reset = 1'd0;
        p23_in = 32'd0;
        p23_write_en = 1'd0;
        p23_clk = 1'd0;
        p23_reset = 1'd0;
        p24_in = 32'd0;
        p24_write_en = 1'd0;
        p24_clk = 1'd0;
        p24_reset = 1'd0;
        p25_in = 32'd0;
        p25_write_en = 1'd0;
        p25_clk = 1'd0;
        p25_reset = 1'd0;
        p26_in = 32'd0;
        p26_write_en = 1'd0;
        p26_clk = 1'd0;
        p26_reset = 1'd0;
        p27_in = 32'd0;
        p27_write_en = 1'd0;
        p27_clk = 1'd0;
        p27_reset = 1'd0;
        p28_in = 32'd0;
        p28_write_en = 1'd0;
        p28_clk = 1'd0;
        p28_reset = 1'd0;
        p29_in = 32'd0;
        p29_write_en = 1'd0;
        p29_clk = 1'd0;
        p29_reset = 1'd0;
        p30_in = 32'd0;
        p30_write_en = 1'd0;
        p30_clk = 1'd0;
        p30_reset = 1'd0;
        p31_in = 32'd0;
        p31_write_en = 1'd0;
        p31_clk = 1'd0;
        p31_reset = 1'd0;
        l0_in = 5'd0;
        l0_write_en = 1'd0;
        l0_clk = 1'd0;
        l0_reset = 1'd0;
        l1_in = 5'd0;
        l1_write_en = 1'd0;
        l1_clk = 1'd0;
        l1_reset = 1'd0;
        l2_in = 5'd0;
        l2_write_en = 1'd0;
        l2_clk = 1'd0;
        l2_reset = 1'd0;
        l3_in = 5'd0;
        l3_write_en = 1'd0;
        l3_clk = 1'd0;
        l3_reset = 1'd0;
        l4_in = 5'd0;
        l4_write_en = 1'd0;
        l4_clk = 1'd0;
        l4_reset = 1'd0;
        l5_in = 5'd0;
        l5_write_en = 1'd0;
        l5_clk = 1'd0;
        l5_reset = 1'd0;
        l6_in = 5'd0;
        l6_write_en = 1'd0;
        l6_clk = 1'd0;
        l6_reset = 1'd0;
        l7_in = 5'd0;
        l7_write_en = 1'd0;
        l7_clk = 1'd0;
        l7_reset = 1'd0;
        l8_in = 5'd0;
        l8_write_en = 1'd0;
        l8_clk = 1'd0;
        l8_reset = 1'd0;
        l9_in = 5'd0;
        l9_write_en = 1'd0;
        l9_clk = 1'd0;
        l9_reset = 1'd0;
        l10_in = 5'd0;
        l10_write_en = 1'd0;
        l10_clk = 1'd0;
        l10_reset = 1'd0;
        l11_in = 5'd0;
        l11_write_en = 1'd0;
        l11_clk = 1'd0;
        l11_reset = 1'd0;
        l12_in = 5'd0;
        l12_write_en = 1'd0;
        l12_clk = 1'd0;
        l12_reset = 1'd0;
        l13_in = 5'd0;
        l13_write_en = 1'd0;
        l13_clk = 1'd0;
        l13_reset = 1'd0;
        l14_in = 5'd0;
        l14_write_en = 1'd0;
        l14_clk = 1'd0;
        l14_reset = 1'd0;
        l15_in = 5'd0;
        l15_write_en = 1'd0;
        l15_clk = 1'd0;
        l15_reset = 1'd0;
        l16_in = 5'd0;
        l16_write_en = 1'd0;
        l16_clk = 1'd0;
        l16_reset = 1'd0;
        l17_in = 5'd0;
        l17_write_en = 1'd0;
        l17_clk = 1'd0;
        l17_reset = 1'd0;
        l18_in = 5'd0;
        l18_write_en = 1'd0;
        l18_clk = 1'd0;
        l18_reset = 1'd0;
        l19_in = 5'd0;
        l19_write_en = 1'd0;
        l19_clk = 1'd0;
        l19_reset = 1'd0;
        l20_in = 5'd0;
        l20_write_en = 1'd0;
        l20_clk = 1'd0;
        l20_reset = 1'd0;
        l21_in = 5'd0;
        l21_write_en = 1'd0;
        l21_clk = 1'd0;
        l21_reset = 1'd0;
        l22_in = 5'd0;
        l22_write_en = 1'd0;
        l22_clk = 1'd0;
        l22_reset = 1'd0;
        l23_in = 5'd0;
        l23_write_en = 1'd0;
        l23_clk = 1'd0;
        l23_reset = 1'd0;
        l24_in = 5'd0;
        l24_write_en = 1'd0;
        l24_clk = 1'd0;
        l24_reset = 1'd0;
        l25_in = 5'd0;
        l25_write_en = 1'd0;
        l25_clk = 1'd0;
        l25_reset = 1'd0;
        l26_in = 5'd0;
        l26_write_en = 1'd0;
        l26_clk = 1'd0;
        l26_reset = 1'd0;
        l27_in = 5'd0;
        l27_write_en = 1'd0;
        l27_clk = 1'd0;
        l27_reset = 1'd0;
        l28_in = 5'd0;
        l28_write_en = 1'd0;
        l28_clk = 1'd0;
        l28_reset = 1'd0;
        l29_in = 5'd0;
        l29_write_en = 1'd0;
        l29_clk = 1'd0;
        l29_reset = 1'd0;
        l30_in = 5'd0;
        l30_write_en = 1'd0;
        l30_clk = 1'd0;
        l30_reset = 1'd0;
        l31_in = 5'd0;
        l31_write_en = 1'd0;
        l31_clk = 1'd0;
        l31_reset = 1'd0;
        is_index0_left = 5'd0;
        is_index0_right = 5'd0;
        is_index1_left = 5'd0;
        is_index1_right = 5'd0;
        is_index2_left = 5'd0;
        is_index2_right = 5'd0;
        is_index3_left = 5'd0;
        is_index3_right = 5'd0;
        is_index4_left = 5'd0;
        is_index4_right = 5'd0;
        is_index5_left = 5'd0;
        is_index5_right = 5'd0;
        is_index6_left = 5'd0;
        is_index6_right = 5'd0;
        is_index7_left = 5'd0;
        is_index7_right = 5'd0;
        is_index8_left = 5'd0;
        is_index8_right = 5'd0;
        is_index9_left = 5'd0;
        is_index9_right = 5'd0;
        is_index10_left = 5'd0;
        is_index10_right = 5'd0;
        is_index11_left = 5'd0;
        is_index11_right = 5'd0;
        is_index12_left = 5'd0;
        is_index12_right = 5'd0;
        is_index13_left = 5'd0;
        is_index13_right = 5'd0;
        is_index14_left = 5'd0;
        is_index14_right = 5'd0;
        is_index15_left = 5'd0;
        is_index15_right = 5'd0;
        is_index16_left = 5'd0;
        is_index16_right = 5'd0;
        is_index17_left = 5'd0;
        is_index17_right = 5'd0;
        is_index18_left = 5'd0;
        is_index18_right = 5'd0;
        is_index19_left = 5'd0;
        is_index19_right = 5'd0;
        is_index20_left = 5'd0;
        is_index20_right = 5'd0;
        is_index21_left = 5'd0;
        is_index21_right = 5'd0;
        is_index22_left = 5'd0;
        is_index22_right = 5'd0;
        is_index23_left = 5'd0;
        is_index23_right = 5'd0;
        is_index24_left = 5'd0;
        is_index24_right = 5'd0;
        is_index25_left = 5'd0;
        is_index25_right = 5'd0;
        is_index26_left = 5'd0;
        is_index26_right = 5'd0;
        is_index27_left = 5'd0;
        is_index27_right = 5'd0;
        is_index28_left = 5'd0;
        is_index28_right = 5'd0;
        is_index29_left = 5'd0;
        is_index29_right = 5'd0;
        is_index30_left = 5'd0;
        is_index30_right = 5'd0;
        is_index31_left = 5'd0;
        is_index31_right = 5'd0;
        zero_index_in = 5'd0;
        zero_index_write_en = 1'd0;
        zero_index_clk = 1'd0;
        zero_index_reset = 1'd0;
        z_eq_left = 6'd0;
        z_eq_right = 6'd0;
        slice_in = 6'd0;
        sub_left = 6'd0;
        sub_right = 6'd0;
        me0_in = 32'd0;
        me0_prefix = 32'd0;
        me0_length = 5'd0;
        me0_go = 1'd0;
        me0_clk = 1'd0;
        me0_reset = 1'd0;
        me1_in = 32'd0;
        me1_prefix = 32'd0;
        me1_length = 5'd0;
        me1_go = 1'd0;
        me1_clk = 1'd0;
        me1_reset = 1'd0;
        me2_in = 32'd0;
        me2_prefix = 32'd0;
        me2_length = 5'd0;
        me2_go = 1'd0;
        me2_clk = 1'd0;
        me2_reset = 1'd0;
        me3_in = 32'd0;
        me3_prefix = 32'd0;
        me3_length = 5'd0;
        me3_go = 1'd0;
        me3_clk = 1'd0;
        me3_reset = 1'd0;
        me4_in = 32'd0;
        me4_prefix = 32'd0;
        me4_length = 5'd0;
        me4_go = 1'd0;
        me4_clk = 1'd0;
        me4_reset = 1'd0;
        me5_in = 32'd0;
        me5_prefix = 32'd0;
        me5_length = 5'd0;
        me5_go = 1'd0;
        me5_clk = 1'd0;
        me5_reset = 1'd0;
        me6_in = 32'd0;
        me6_prefix = 32'd0;
        me6_length = 5'd0;
        me6_go = 1'd0;
        me6_clk = 1'd0;
        me6_reset = 1'd0;
        me7_in = 32'd0;
        me7_prefix = 32'd0;
        me7_length = 5'd0;
        me7_go = 1'd0;
        me7_clk = 1'd0;
        me7_reset = 1'd0;
        me8_in = 32'd0;
        me8_prefix = 32'd0;
        me8_length = 5'd0;
        me8_go = 1'd0;
        me8_clk = 1'd0;
        me8_reset = 1'd0;
        me9_in = 32'd0;
        me9_prefix = 32'd0;
        me9_length = 5'd0;
        me9_go = 1'd0;
        me9_clk = 1'd0;
        me9_reset = 1'd0;
        me10_in = 32'd0;
        me10_prefix = 32'd0;
        me10_length = 5'd0;
        me10_go = 1'd0;
        me10_clk = 1'd0;
        me10_reset = 1'd0;
        me11_in = 32'd0;
        me11_prefix = 32'd0;
        me11_length = 5'd0;
        me11_go = 1'd0;
        me11_clk = 1'd0;
        me11_reset = 1'd0;
        me12_in = 32'd0;
        me12_prefix = 32'd0;
        me12_length = 5'd0;
        me12_go = 1'd0;
        me12_clk = 1'd0;
        me12_reset = 1'd0;
        me13_in = 32'd0;
        me13_prefix = 32'd0;
        me13_length = 5'd0;
        me13_go = 1'd0;
        me13_clk = 1'd0;
        me13_reset = 1'd0;
        me14_in = 32'd0;
        me14_prefix = 32'd0;
        me14_length = 5'd0;
        me14_go = 1'd0;
        me14_clk = 1'd0;
        me14_reset = 1'd0;
        me15_in = 32'd0;
        me15_prefix = 32'd0;
        me15_length = 5'd0;
        me15_go = 1'd0;
        me15_clk = 1'd0;
        me15_reset = 1'd0;
        me16_in = 32'd0;
        me16_prefix = 32'd0;
        me16_length = 5'd0;
        me16_go = 1'd0;
        me16_clk = 1'd0;
        me16_reset = 1'd0;
        me17_in = 32'd0;
        me17_prefix = 32'd0;
        me17_length = 5'd0;
        me17_go = 1'd0;
        me17_clk = 1'd0;
        me17_reset = 1'd0;
        me18_in = 32'd0;
        me18_prefix = 32'd0;
        me18_length = 5'd0;
        me18_go = 1'd0;
        me18_clk = 1'd0;
        me18_reset = 1'd0;
        me19_in = 32'd0;
        me19_prefix = 32'd0;
        me19_length = 5'd0;
        me19_go = 1'd0;
        me19_clk = 1'd0;
        me19_reset = 1'd0;
        me20_in = 32'd0;
        me20_prefix = 32'd0;
        me20_length = 5'd0;
        me20_go = 1'd0;
        me20_clk = 1'd0;
        me20_reset = 1'd0;
        me21_in = 32'd0;
        me21_prefix = 32'd0;
        me21_length = 5'd0;
        me21_go = 1'd0;
        me21_clk = 1'd0;
        me21_reset = 1'd0;
        me22_in = 32'd0;
        me22_prefix = 32'd0;
        me22_length = 5'd0;
        me22_go = 1'd0;
        me22_clk = 1'd0;
        me22_reset = 1'd0;
        me23_in = 32'd0;
        me23_prefix = 32'd0;
        me23_length = 5'd0;
        me23_go = 1'd0;
        me23_clk = 1'd0;
        me23_reset = 1'd0;
        me24_in = 32'd0;
        me24_prefix = 32'd0;
        me24_length = 5'd0;
        me24_go = 1'd0;
        me24_clk = 1'd0;
        me24_reset = 1'd0;
        me25_in = 32'd0;
        me25_prefix = 32'd0;
        me25_length = 5'd0;
        me25_go = 1'd0;
        me25_clk = 1'd0;
        me25_reset = 1'd0;
        me26_in = 32'd0;
        me26_prefix = 32'd0;
        me26_length = 5'd0;
        me26_go = 1'd0;
        me26_clk = 1'd0;
        me26_reset = 1'd0;
        me27_in = 32'd0;
        me27_prefix = 32'd0;
        me27_length = 5'd0;
        me27_go = 1'd0;
        me27_clk = 1'd0;
        me27_reset = 1'd0;
        me28_in = 32'd0;
        me28_prefix = 32'd0;
        me28_length = 5'd0;
        me28_go = 1'd0;
        me28_clk = 1'd0;
        me28_reset = 1'd0;
        me29_in = 32'd0;
        me29_prefix = 32'd0;
        me29_length = 5'd0;
        me29_go = 1'd0;
        me29_clk = 1'd0;
        me29_reset = 1'd0;
        me30_in = 32'd0;
        me30_prefix = 32'd0;
        me30_length = 5'd0;
        me30_go = 1'd0;
        me30_clk = 1'd0;
        me30_reset = 1'd0;
        me31_in = 32'd0;
        me31_prefix = 32'd0;
        me31_length = 5'd0;
        me31_go = 1'd0;
        me31_clk = 1'd0;
        me31_reset = 1'd0;
        ce00_lenA = 5'd0;
        ce00_lenB = 5'd0;
        ce00_addrA = 5'd0;
        ce00_addrB = 5'd0;
        ce00_mlA = 1'd0;
        ce00_mlB = 1'd0;
        ce00_go = 1'd0;
        ce00_clk = 1'd0;
        ce00_reset = 1'd0;
        ce01_lenA = 5'd0;
        ce01_lenB = 5'd0;
        ce01_addrA = 5'd0;
        ce01_addrB = 5'd0;
        ce01_mlA = 1'd0;
        ce01_mlB = 1'd0;
        ce01_go = 1'd0;
        ce01_clk = 1'd0;
        ce01_reset = 1'd0;
        ce02_lenA = 5'd0;
        ce02_lenB = 5'd0;
        ce02_addrA = 5'd0;
        ce02_addrB = 5'd0;
        ce02_mlA = 1'd0;
        ce02_mlB = 1'd0;
        ce02_go = 1'd0;
        ce02_clk = 1'd0;
        ce02_reset = 1'd0;
        ce03_lenA = 5'd0;
        ce03_lenB = 5'd0;
        ce03_addrA = 5'd0;
        ce03_addrB = 5'd0;
        ce03_mlA = 1'd0;
        ce03_mlB = 1'd0;
        ce03_go = 1'd0;
        ce03_clk = 1'd0;
        ce03_reset = 1'd0;
        ce04_lenA = 5'd0;
        ce04_lenB = 5'd0;
        ce04_addrA = 5'd0;
        ce04_addrB = 5'd0;
        ce04_mlA = 1'd0;
        ce04_mlB = 1'd0;
        ce04_go = 1'd0;
        ce04_clk = 1'd0;
        ce04_reset = 1'd0;
        ce05_lenA = 5'd0;
        ce05_lenB = 5'd0;
        ce05_addrA = 5'd0;
        ce05_addrB = 5'd0;
        ce05_mlA = 1'd0;
        ce05_mlB = 1'd0;
        ce05_go = 1'd0;
        ce05_clk = 1'd0;
        ce05_reset = 1'd0;
        ce06_lenA = 5'd0;
        ce06_lenB = 5'd0;
        ce06_addrA = 5'd0;
        ce06_addrB = 5'd0;
        ce06_mlA = 1'd0;
        ce06_mlB = 1'd0;
        ce06_go = 1'd0;
        ce06_clk = 1'd0;
        ce06_reset = 1'd0;
        ce07_lenA = 5'd0;
        ce07_lenB = 5'd0;
        ce07_addrA = 5'd0;
        ce07_addrB = 5'd0;
        ce07_mlA = 1'd0;
        ce07_mlB = 1'd0;
        ce07_go = 1'd0;
        ce07_clk = 1'd0;
        ce07_reset = 1'd0;
        ce08_lenA = 5'd0;
        ce08_lenB = 5'd0;
        ce08_addrA = 5'd0;
        ce08_addrB = 5'd0;
        ce08_mlA = 1'd0;
        ce08_mlB = 1'd0;
        ce08_go = 1'd0;
        ce08_clk = 1'd0;
        ce08_reset = 1'd0;
        ce09_lenA = 5'd0;
        ce09_lenB = 5'd0;
        ce09_addrA = 5'd0;
        ce09_addrB = 5'd0;
        ce09_mlA = 1'd0;
        ce09_mlB = 1'd0;
        ce09_go = 1'd0;
        ce09_clk = 1'd0;
        ce09_reset = 1'd0;
        ce010_lenA = 5'd0;
        ce010_lenB = 5'd0;
        ce010_addrA = 5'd0;
        ce010_addrB = 5'd0;
        ce010_mlA = 1'd0;
        ce010_mlB = 1'd0;
        ce010_go = 1'd0;
        ce010_clk = 1'd0;
        ce010_reset = 1'd0;
        ce011_lenA = 5'd0;
        ce011_lenB = 5'd0;
        ce011_addrA = 5'd0;
        ce011_addrB = 5'd0;
        ce011_mlA = 1'd0;
        ce011_mlB = 1'd0;
        ce011_go = 1'd0;
        ce011_clk = 1'd0;
        ce011_reset = 1'd0;
        ce012_lenA = 5'd0;
        ce012_lenB = 5'd0;
        ce012_addrA = 5'd0;
        ce012_addrB = 5'd0;
        ce012_mlA = 1'd0;
        ce012_mlB = 1'd0;
        ce012_go = 1'd0;
        ce012_clk = 1'd0;
        ce012_reset = 1'd0;
        ce013_lenA = 5'd0;
        ce013_lenB = 5'd0;
        ce013_addrA = 5'd0;
        ce013_addrB = 5'd0;
        ce013_mlA = 1'd0;
        ce013_mlB = 1'd0;
        ce013_go = 1'd0;
        ce013_clk = 1'd0;
        ce013_reset = 1'd0;
        ce014_lenA = 5'd0;
        ce014_lenB = 5'd0;
        ce014_addrA = 5'd0;
        ce014_addrB = 5'd0;
        ce014_mlA = 1'd0;
        ce014_mlB = 1'd0;
        ce014_go = 1'd0;
        ce014_clk = 1'd0;
        ce014_reset = 1'd0;
        ce015_lenA = 5'd0;
        ce015_lenB = 5'd0;
        ce015_addrA = 5'd0;
        ce015_addrB = 5'd0;
        ce015_mlA = 1'd0;
        ce015_mlB = 1'd0;
        ce015_go = 1'd0;
        ce015_clk = 1'd0;
        ce015_reset = 1'd0;
        ce10_lenA = 5'd0;
        ce10_lenB = 5'd0;
        ce10_addrA = 5'd0;
        ce10_addrB = 5'd0;
        ce10_mlA = 1'd0;
        ce10_mlB = 1'd0;
        ce10_go = 1'd0;
        ce10_clk = 1'd0;
        ce10_reset = 1'd0;
        ce11_lenA = 5'd0;
        ce11_lenB = 5'd0;
        ce11_addrA = 5'd0;
        ce11_addrB = 5'd0;
        ce11_mlA = 1'd0;
        ce11_mlB = 1'd0;
        ce11_go = 1'd0;
        ce11_clk = 1'd0;
        ce11_reset = 1'd0;
        ce12_lenA = 5'd0;
        ce12_lenB = 5'd0;
        ce12_addrA = 5'd0;
        ce12_addrB = 5'd0;
        ce12_mlA = 1'd0;
        ce12_mlB = 1'd0;
        ce12_go = 1'd0;
        ce12_clk = 1'd0;
        ce12_reset = 1'd0;
        ce13_lenA = 5'd0;
        ce13_lenB = 5'd0;
        ce13_addrA = 5'd0;
        ce13_addrB = 5'd0;
        ce13_mlA = 1'd0;
        ce13_mlB = 1'd0;
        ce13_go = 1'd0;
        ce13_clk = 1'd0;
        ce13_reset = 1'd0;
        ce14_lenA = 5'd0;
        ce14_lenB = 5'd0;
        ce14_addrA = 5'd0;
        ce14_addrB = 5'd0;
        ce14_mlA = 1'd0;
        ce14_mlB = 1'd0;
        ce14_go = 1'd0;
        ce14_clk = 1'd0;
        ce14_reset = 1'd0;
        ce15_lenA = 5'd0;
        ce15_lenB = 5'd0;
        ce15_addrA = 5'd0;
        ce15_addrB = 5'd0;
        ce15_mlA = 1'd0;
        ce15_mlB = 1'd0;
        ce15_go = 1'd0;
        ce15_clk = 1'd0;
        ce15_reset = 1'd0;
        ce16_lenA = 5'd0;
        ce16_lenB = 5'd0;
        ce16_addrA = 5'd0;
        ce16_addrB = 5'd0;
        ce16_mlA = 1'd0;
        ce16_mlB = 1'd0;
        ce16_go = 1'd0;
        ce16_clk = 1'd0;
        ce16_reset = 1'd0;
        ce17_lenA = 5'd0;
        ce17_lenB = 5'd0;
        ce17_addrA = 5'd0;
        ce17_addrB = 5'd0;
        ce17_mlA = 1'd0;
        ce17_mlB = 1'd0;
        ce17_go = 1'd0;
        ce17_clk = 1'd0;
        ce17_reset = 1'd0;
        ce20_lenA = 5'd0;
        ce20_lenB = 5'd0;
        ce20_addrA = 5'd0;
        ce20_addrB = 5'd0;
        ce20_mlA = 1'd0;
        ce20_mlB = 1'd0;
        ce20_go = 1'd0;
        ce20_clk = 1'd0;
        ce20_reset = 1'd0;
        ce21_lenA = 5'd0;
        ce21_lenB = 5'd0;
        ce21_addrA = 5'd0;
        ce21_addrB = 5'd0;
        ce21_mlA = 1'd0;
        ce21_mlB = 1'd0;
        ce21_go = 1'd0;
        ce21_clk = 1'd0;
        ce21_reset = 1'd0;
        ce22_lenA = 5'd0;
        ce22_lenB = 5'd0;
        ce22_addrA = 5'd0;
        ce22_addrB = 5'd0;
        ce22_mlA = 1'd0;
        ce22_mlB = 1'd0;
        ce22_go = 1'd0;
        ce22_clk = 1'd0;
        ce22_reset = 1'd0;
        ce23_lenA = 5'd0;
        ce23_lenB = 5'd0;
        ce23_addrA = 5'd0;
        ce23_addrB = 5'd0;
        ce23_mlA = 1'd0;
        ce23_mlB = 1'd0;
        ce23_go = 1'd0;
        ce23_clk = 1'd0;
        ce23_reset = 1'd0;
        ce30_lenA = 5'd0;
        ce30_lenB = 5'd0;
        ce30_addrA = 5'd0;
        ce30_addrB = 5'd0;
        ce30_mlA = 1'd0;
        ce30_mlB = 1'd0;
        ce30_go = 1'd0;
        ce30_clk = 1'd0;
        ce30_reset = 1'd0;
        ce31_lenA = 5'd0;
        ce31_lenB = 5'd0;
        ce31_addrA = 5'd0;
        ce31_addrB = 5'd0;
        ce31_mlA = 1'd0;
        ce31_mlB = 1'd0;
        ce31_go = 1'd0;
        ce31_clk = 1'd0;
        ce31_reset = 1'd0;
        ce40_lenA = 5'd0;
        ce40_lenB = 5'd0;
        ce40_addrA = 5'd0;
        ce40_addrB = 5'd0;
        ce40_mlA = 1'd0;
        ce40_mlB = 1'd0;
        ce40_go = 1'd0;
        ce40_clk = 1'd0;
        ce40_reset = 1'd0;
        comb_reg0_in = 1'd0;
        comb_reg0_write_en = 1'd0;
        comb_reg0_clk = 1'd0;
        comb_reg0_reset = 1'd0;
        comb_reg1_in = 1'd0;
        comb_reg1_write_en = 1'd0;
        comb_reg1_clk = 1'd0;
        comb_reg1_reset = 1'd0;
        comb_reg2_in = 1'd0;
        comb_reg2_write_en = 1'd0;
        comb_reg2_clk = 1'd0;
        comb_reg2_reset = 1'd0;
        comb_reg3_in = 1'd0;
        comb_reg3_write_en = 1'd0;
        comb_reg3_clk = 1'd0;
        comb_reg3_reset = 1'd0;
        comb_reg4_in = 1'd0;
        comb_reg4_write_en = 1'd0;
        comb_reg4_clk = 1'd0;
        comb_reg4_reset = 1'd0;
        comb_reg5_in = 1'd0;
        comb_reg5_write_en = 1'd0;
        comb_reg5_clk = 1'd0;
        comb_reg5_reset = 1'd0;
        comb_reg6_in = 1'd0;
        comb_reg6_write_en = 1'd0;
        comb_reg6_clk = 1'd0;
        comb_reg6_reset = 1'd0;
        comb_reg7_in = 1'd0;
        comb_reg7_write_en = 1'd0;
        comb_reg7_clk = 1'd0;
        comb_reg7_reset = 1'd0;
        comb_reg8_in = 1'd0;
        comb_reg8_write_en = 1'd0;
        comb_reg8_clk = 1'd0;
        comb_reg8_reset = 1'd0;
        comb_reg9_in = 1'd0;
        comb_reg9_write_en = 1'd0;
        comb_reg9_clk = 1'd0;
        comb_reg9_reset = 1'd0;
        comb_reg10_in = 1'd0;
        comb_reg10_write_en = 1'd0;
        comb_reg10_clk = 1'd0;
        comb_reg10_reset = 1'd0;
        comb_reg11_in = 1'd0;
        comb_reg11_write_en = 1'd0;
        comb_reg11_clk = 1'd0;
        comb_reg11_reset = 1'd0;
        comb_reg12_in = 1'd0;
        comb_reg12_write_en = 1'd0;
        comb_reg12_clk = 1'd0;
        comb_reg12_reset = 1'd0;
        comb_reg13_in = 1'd0;
        comb_reg13_write_en = 1'd0;
        comb_reg13_clk = 1'd0;
        comb_reg13_reset = 1'd0;
        comb_reg14_in = 1'd0;
        comb_reg14_write_en = 1'd0;
        comb_reg14_clk = 1'd0;
        comb_reg14_reset = 1'd0;
        comb_reg15_in = 1'd0;
        comb_reg15_write_en = 1'd0;
        comb_reg15_clk = 1'd0;
        comb_reg15_reset = 1'd0;
        comb_reg16_in = 1'd0;
        comb_reg16_write_en = 1'd0;
        comb_reg16_clk = 1'd0;
        comb_reg16_reset = 1'd0;
        comb_reg17_in = 1'd0;
        comb_reg17_write_en = 1'd0;
        comb_reg17_clk = 1'd0;
        comb_reg17_reset = 1'd0;
        comb_reg18_in = 1'd0;
        comb_reg18_write_en = 1'd0;
        comb_reg18_clk = 1'd0;
        comb_reg18_reset = 1'd0;
        comb_reg19_in = 1'd0;
        comb_reg19_write_en = 1'd0;
        comb_reg19_clk = 1'd0;
        comb_reg19_reset = 1'd0;
        comb_reg20_in = 1'd0;
        comb_reg20_write_en = 1'd0;
        comb_reg20_clk = 1'd0;
        comb_reg20_reset = 1'd0;
        comb_reg21_in = 1'd0;
        comb_reg21_write_en = 1'd0;
        comb_reg21_clk = 1'd0;
        comb_reg21_reset = 1'd0;
        comb_reg22_in = 1'd0;
        comb_reg22_write_en = 1'd0;
        comb_reg22_clk = 1'd0;
        comb_reg22_reset = 1'd0;
        comb_reg23_in = 1'd0;
        comb_reg23_write_en = 1'd0;
        comb_reg23_clk = 1'd0;
        comb_reg23_reset = 1'd0;
        comb_reg24_in = 1'd0;
        comb_reg24_write_en = 1'd0;
        comb_reg24_clk = 1'd0;
        comb_reg24_reset = 1'd0;
        comb_reg25_in = 1'd0;
        comb_reg25_write_en = 1'd0;
        comb_reg25_clk = 1'd0;
        comb_reg25_reset = 1'd0;
        comb_reg26_in = 1'd0;
        comb_reg26_write_en = 1'd0;
        comb_reg26_clk = 1'd0;
        comb_reg26_reset = 1'd0;
        comb_reg27_in = 1'd0;
        comb_reg27_write_en = 1'd0;
        comb_reg27_clk = 1'd0;
        comb_reg27_reset = 1'd0;
        comb_reg28_in = 1'd0;
        comb_reg28_write_en = 1'd0;
        comb_reg28_clk = 1'd0;
        comb_reg28_reset = 1'd0;
        comb_reg29_in = 1'd0;
        comb_reg29_write_en = 1'd0;
        comb_reg29_clk = 1'd0;
        comb_reg29_reset = 1'd0;
        comb_reg30_in = 1'd0;
        comb_reg30_write_en = 1'd0;
        comb_reg30_clk = 1'd0;
        comb_reg30_reset = 1'd0;
        comb_reg31_in = 1'd0;
        comb_reg31_write_en = 1'd0;
        comb_reg31_clk = 1'd0;
        comb_reg31_reset = 1'd0;
        out_in = 5'd0;
        out_write_en = 1'd0;
        out_clk = 1'd0;
        out_reset = 1'd0;
        fsm_in = 2'd0;
        fsm_write_en = 1'd0;
        fsm_clk = 1'd0;
        fsm_reset = 1'd0;
        pd_in = 1'd0;
        pd_write_en = 1'd0;
        pd_clk = 1'd0;
        pd_reset = 1'd0;
        fsm0_in = 2'd0;
        fsm0_write_en = 1'd0;
        fsm0_clk = 1'd0;
        fsm0_reset = 1'd0;
        pd0_in = 1'd0;
        pd0_write_en = 1'd0;
        pd0_clk = 1'd0;
        pd0_reset = 1'd0;
        fsm1_in = 2'd0;
        fsm1_write_en = 1'd0;
        fsm1_clk = 1'd0;
        fsm1_reset = 1'd0;
        pd1_in = 1'd0;
        pd1_write_en = 1'd0;
        pd1_clk = 1'd0;
        pd1_reset = 1'd0;
        fsm2_in = 2'd0;
        fsm2_write_en = 1'd0;
        fsm2_clk = 1'd0;
        fsm2_reset = 1'd0;
        pd2_in = 1'd0;
        pd2_write_en = 1'd0;
        pd2_clk = 1'd0;
        pd2_reset = 1'd0;
        fsm3_in = 2'd0;
        fsm3_write_en = 1'd0;
        fsm3_clk = 1'd0;
        fsm3_reset = 1'd0;
        pd3_in = 1'd0;
        pd3_write_en = 1'd0;
        pd3_clk = 1'd0;
        pd3_reset = 1'd0;
        fsm4_in = 2'd0;
        fsm4_write_en = 1'd0;
        fsm4_clk = 1'd0;
        fsm4_reset = 1'd0;
        pd4_in = 1'd0;
        pd4_write_en = 1'd0;
        pd4_clk = 1'd0;
        pd4_reset = 1'd0;
        fsm5_in = 2'd0;
        fsm5_write_en = 1'd0;
        fsm5_clk = 1'd0;
        fsm5_reset = 1'd0;
        pd5_in = 1'd0;
        pd5_write_en = 1'd0;
        pd5_clk = 1'd0;
        pd5_reset = 1'd0;
        fsm6_in = 2'd0;
        fsm6_write_en = 1'd0;
        fsm6_clk = 1'd0;
        fsm6_reset = 1'd0;
        pd6_in = 1'd0;
        pd6_write_en = 1'd0;
        pd6_clk = 1'd0;
        pd6_reset = 1'd0;
        fsm7_in = 2'd0;
        fsm7_write_en = 1'd0;
        fsm7_clk = 1'd0;
        fsm7_reset = 1'd0;
        pd7_in = 1'd0;
        pd7_write_en = 1'd0;
        pd7_clk = 1'd0;
        pd7_reset = 1'd0;
        fsm8_in = 2'd0;
        fsm8_write_en = 1'd0;
        fsm8_clk = 1'd0;
        fsm8_reset = 1'd0;
        pd8_in = 1'd0;
        pd8_write_en = 1'd0;
        pd8_clk = 1'd0;
        pd8_reset = 1'd0;
        fsm9_in = 2'd0;
        fsm9_write_en = 1'd0;
        fsm9_clk = 1'd0;
        fsm9_reset = 1'd0;
        pd9_in = 1'd0;
        pd9_write_en = 1'd0;
        pd9_clk = 1'd0;
        pd9_reset = 1'd0;
        fsm10_in = 2'd0;
        fsm10_write_en = 1'd0;
        fsm10_clk = 1'd0;
        fsm10_reset = 1'd0;
        pd10_in = 1'd0;
        pd10_write_en = 1'd0;
        pd10_clk = 1'd0;
        pd10_reset = 1'd0;
        fsm11_in = 2'd0;
        fsm11_write_en = 1'd0;
        fsm11_clk = 1'd0;
        fsm11_reset = 1'd0;
        pd11_in = 1'd0;
        pd11_write_en = 1'd0;
        pd11_clk = 1'd0;
        pd11_reset = 1'd0;
        fsm12_in = 2'd0;
        fsm12_write_en = 1'd0;
        fsm12_clk = 1'd0;
        fsm12_reset = 1'd0;
        pd12_in = 1'd0;
        pd12_write_en = 1'd0;
        pd12_clk = 1'd0;
        pd12_reset = 1'd0;
        fsm13_in = 2'd0;
        fsm13_write_en = 1'd0;
        fsm13_clk = 1'd0;
        fsm13_reset = 1'd0;
        pd13_in = 1'd0;
        pd13_write_en = 1'd0;
        pd13_clk = 1'd0;
        pd13_reset = 1'd0;
        fsm14_in = 2'd0;
        fsm14_write_en = 1'd0;
        fsm14_clk = 1'd0;
        fsm14_reset = 1'd0;
        pd14_in = 1'd0;
        pd14_write_en = 1'd0;
        pd14_clk = 1'd0;
        pd14_reset = 1'd0;
        fsm15_in = 2'd0;
        fsm15_write_en = 1'd0;
        fsm15_clk = 1'd0;
        fsm15_reset = 1'd0;
        pd15_in = 1'd0;
        pd15_write_en = 1'd0;
        pd15_clk = 1'd0;
        pd15_reset = 1'd0;
        fsm16_in = 2'd0;
        fsm16_write_en = 1'd0;
        fsm16_clk = 1'd0;
        fsm16_reset = 1'd0;
        pd16_in = 1'd0;
        pd16_write_en = 1'd0;
        pd16_clk = 1'd0;
        pd16_reset = 1'd0;
        fsm17_in = 2'd0;
        fsm17_write_en = 1'd0;
        fsm17_clk = 1'd0;
        fsm17_reset = 1'd0;
        pd17_in = 1'd0;
        pd17_write_en = 1'd0;
        pd17_clk = 1'd0;
        pd17_reset = 1'd0;
        fsm18_in = 2'd0;
        fsm18_write_en = 1'd0;
        fsm18_clk = 1'd0;
        fsm18_reset = 1'd0;
        pd18_in = 1'd0;
        pd18_write_en = 1'd0;
        pd18_clk = 1'd0;
        pd18_reset = 1'd0;
        fsm19_in = 2'd0;
        fsm19_write_en = 1'd0;
        fsm19_clk = 1'd0;
        fsm19_reset = 1'd0;
        pd19_in = 1'd0;
        pd19_write_en = 1'd0;
        pd19_clk = 1'd0;
        pd19_reset = 1'd0;
        fsm20_in = 2'd0;
        fsm20_write_en = 1'd0;
        fsm20_clk = 1'd0;
        fsm20_reset = 1'd0;
        pd20_in = 1'd0;
        pd20_write_en = 1'd0;
        pd20_clk = 1'd0;
        pd20_reset = 1'd0;
        fsm21_in = 2'd0;
        fsm21_write_en = 1'd0;
        fsm21_clk = 1'd0;
        fsm21_reset = 1'd0;
        pd21_in = 1'd0;
        pd21_write_en = 1'd0;
        pd21_clk = 1'd0;
        pd21_reset = 1'd0;
        fsm22_in = 2'd0;
        fsm22_write_en = 1'd0;
        fsm22_clk = 1'd0;
        fsm22_reset = 1'd0;
        pd22_in = 1'd0;
        pd22_write_en = 1'd0;
        pd22_clk = 1'd0;
        pd22_reset = 1'd0;
        fsm23_in = 2'd0;
        fsm23_write_en = 1'd0;
        fsm23_clk = 1'd0;
        fsm23_reset = 1'd0;
        pd23_in = 1'd0;
        pd23_write_en = 1'd0;
        pd23_clk = 1'd0;
        pd23_reset = 1'd0;
        fsm24_in = 2'd0;
        fsm24_write_en = 1'd0;
        fsm24_clk = 1'd0;
        fsm24_reset = 1'd0;
        pd24_in = 1'd0;
        pd24_write_en = 1'd0;
        pd24_clk = 1'd0;
        pd24_reset = 1'd0;
        fsm25_in = 2'd0;
        fsm25_write_en = 1'd0;
        fsm25_clk = 1'd0;
        fsm25_reset = 1'd0;
        pd25_in = 1'd0;
        pd25_write_en = 1'd0;
        pd25_clk = 1'd0;
        pd25_reset = 1'd0;
        fsm26_in = 2'd0;
        fsm26_write_en = 1'd0;
        fsm26_clk = 1'd0;
        fsm26_reset = 1'd0;
        pd26_in = 1'd0;
        pd26_write_en = 1'd0;
        pd26_clk = 1'd0;
        pd26_reset = 1'd0;
        fsm27_in = 2'd0;
        fsm27_write_en = 1'd0;
        fsm27_clk = 1'd0;
        fsm27_reset = 1'd0;
        pd27_in = 1'd0;
        pd27_write_en = 1'd0;
        pd27_clk = 1'd0;
        pd27_reset = 1'd0;
        fsm28_in = 2'd0;
        fsm28_write_en = 1'd0;
        fsm28_clk = 1'd0;
        fsm28_reset = 1'd0;
        pd28_in = 1'd0;
        pd28_write_en = 1'd0;
        pd28_clk = 1'd0;
        pd28_reset = 1'd0;
        fsm29_in = 2'd0;
        fsm29_write_en = 1'd0;
        fsm29_clk = 1'd0;
        fsm29_reset = 1'd0;
        pd29_in = 1'd0;
        pd29_write_en = 1'd0;
        pd29_clk = 1'd0;
        pd29_reset = 1'd0;
        fsm30_in = 2'd0;
        fsm30_write_en = 1'd0;
        fsm30_clk = 1'd0;
        fsm30_reset = 1'd0;
        pd30_in = 1'd0;
        pd30_write_en = 1'd0;
        pd30_clk = 1'd0;
        pd30_reset = 1'd0;
        pd31_in = 1'd0;
        pd31_write_en = 1'd0;
        pd31_clk = 1'd0;
        pd31_reset = 1'd0;
        pd32_in = 1'd0;
        pd32_write_en = 1'd0;
        pd32_clk = 1'd0;
        pd32_reset = 1'd0;
        pd33_in = 1'd0;
        pd33_write_en = 1'd0;
        pd33_clk = 1'd0;
        pd33_reset = 1'd0;
        pd34_in = 1'd0;
        pd34_write_en = 1'd0;
        pd34_clk = 1'd0;
        pd34_reset = 1'd0;
        pd35_in = 1'd0;
        pd35_write_en = 1'd0;
        pd35_clk = 1'd0;
        pd35_reset = 1'd0;
        pd36_in = 1'd0;
        pd36_write_en = 1'd0;
        pd36_clk = 1'd0;
        pd36_reset = 1'd0;
        pd37_in = 1'd0;
        pd37_write_en = 1'd0;
        pd37_clk = 1'd0;
        pd37_reset = 1'd0;
        pd38_in = 1'd0;
        pd38_write_en = 1'd0;
        pd38_clk = 1'd0;
        pd38_reset = 1'd0;
        pd39_in = 1'd0;
        pd39_write_en = 1'd0;
        pd39_clk = 1'd0;
        pd39_reset = 1'd0;
        pd40_in = 1'd0;
        pd40_write_en = 1'd0;
        pd40_clk = 1'd0;
        pd40_reset = 1'd0;
        pd41_in = 1'd0;
        pd41_write_en = 1'd0;
        pd41_clk = 1'd0;
        pd41_reset = 1'd0;
        pd42_in = 1'd0;
        pd42_write_en = 1'd0;
        pd42_clk = 1'd0;
        pd42_reset = 1'd0;
        pd43_in = 1'd0;
        pd43_write_en = 1'd0;
        pd43_clk = 1'd0;
        pd43_reset = 1'd0;
        pd44_in = 1'd0;
        pd44_write_en = 1'd0;
        pd44_clk = 1'd0;
        pd44_reset = 1'd0;
        pd45_in = 1'd0;
        pd45_write_en = 1'd0;
        pd45_clk = 1'd0;
        pd45_reset = 1'd0;
        pd46_in = 1'd0;
        pd46_write_en = 1'd0;
        pd46_clk = 1'd0;
        pd46_reset = 1'd0;
        pd47_in = 1'd0;
        pd47_write_en = 1'd0;
        pd47_clk = 1'd0;
        pd47_reset = 1'd0;
        pd48_in = 1'd0;
        pd48_write_en = 1'd0;
        pd48_clk = 1'd0;
        pd48_reset = 1'd0;
        pd49_in = 1'd0;
        pd49_write_en = 1'd0;
        pd49_clk = 1'd0;
        pd49_reset = 1'd0;
        pd50_in = 1'd0;
        pd50_write_en = 1'd0;
        pd50_clk = 1'd0;
        pd50_reset = 1'd0;
        pd51_in = 1'd0;
        pd51_write_en = 1'd0;
        pd51_clk = 1'd0;
        pd51_reset = 1'd0;
        pd52_in = 1'd0;
        pd52_write_en = 1'd0;
        pd52_clk = 1'd0;
        pd52_reset = 1'd0;
        pd53_in = 1'd0;
        pd53_write_en = 1'd0;
        pd53_clk = 1'd0;
        pd53_reset = 1'd0;
        pd54_in = 1'd0;
        pd54_write_en = 1'd0;
        pd54_clk = 1'd0;
        pd54_reset = 1'd0;
        pd55_in = 1'd0;
        pd55_write_en = 1'd0;
        pd55_clk = 1'd0;
        pd55_reset = 1'd0;
        pd56_in = 1'd0;
        pd56_write_en = 1'd0;
        pd56_clk = 1'd0;
        pd56_reset = 1'd0;
        pd57_in = 1'd0;
        pd57_write_en = 1'd0;
        pd57_clk = 1'd0;
        pd57_reset = 1'd0;
        pd58_in = 1'd0;
        pd58_write_en = 1'd0;
        pd58_clk = 1'd0;
        pd58_reset = 1'd0;
        pd59_in = 1'd0;
        pd59_write_en = 1'd0;
        pd59_clk = 1'd0;
        pd59_reset = 1'd0;
        pd60_in = 1'd0;
        pd60_write_en = 1'd0;
        pd60_clk = 1'd0;
        pd60_reset = 1'd0;
        pd61_in = 1'd0;
        pd61_write_en = 1'd0;
        pd61_clk = 1'd0;
        pd61_reset = 1'd0;
        pd62_in = 1'd0;
        pd62_write_en = 1'd0;
        pd62_clk = 1'd0;
        pd62_reset = 1'd0;
        pd63_in = 1'd0;
        pd63_write_en = 1'd0;
        pd63_clk = 1'd0;
        pd63_reset = 1'd0;
        pd64_in = 1'd0;
        pd64_write_en = 1'd0;
        pd64_clk = 1'd0;
        pd64_reset = 1'd0;
        pd65_in = 1'd0;
        pd65_write_en = 1'd0;
        pd65_clk = 1'd0;
        pd65_reset = 1'd0;
        pd66_in = 1'd0;
        pd66_write_en = 1'd0;
        pd66_clk = 1'd0;
        pd66_reset = 1'd0;
        pd67_in = 1'd0;
        pd67_write_en = 1'd0;
        pd67_clk = 1'd0;
        pd67_reset = 1'd0;
        pd68_in = 1'd0;
        pd68_write_en = 1'd0;
        pd68_clk = 1'd0;
        pd68_reset = 1'd0;
        pd69_in = 1'd0;
        pd69_write_en = 1'd0;
        pd69_clk = 1'd0;
        pd69_reset = 1'd0;
        pd70_in = 1'd0;
        pd70_write_en = 1'd0;
        pd70_clk = 1'd0;
        pd70_reset = 1'd0;
        pd71_in = 1'd0;
        pd71_write_en = 1'd0;
        pd71_clk = 1'd0;
        pd71_reset = 1'd0;
        pd72_in = 1'd0;
        pd72_write_en = 1'd0;
        pd72_clk = 1'd0;
        pd72_reset = 1'd0;
        pd73_in = 1'd0;
        pd73_write_en = 1'd0;
        pd73_clk = 1'd0;
        pd73_reset = 1'd0;
        pd74_in = 1'd0;
        pd74_write_en = 1'd0;
        pd74_clk = 1'd0;
        pd74_reset = 1'd0;
        pd75_in = 1'd0;
        pd75_write_en = 1'd0;
        pd75_clk = 1'd0;
        pd75_reset = 1'd0;
        pd76_in = 1'd0;
        pd76_write_en = 1'd0;
        pd76_clk = 1'd0;
        pd76_reset = 1'd0;
        pd77_in = 1'd0;
        pd77_write_en = 1'd0;
        pd77_clk = 1'd0;
        pd77_reset = 1'd0;
        pd78_in = 1'd0;
        pd78_write_en = 1'd0;
        pd78_clk = 1'd0;
        pd78_reset = 1'd0;
        pd79_in = 1'd0;
        pd79_write_en = 1'd0;
        pd79_clk = 1'd0;
        pd79_reset = 1'd0;
        pd80_in = 1'd0;
        pd80_write_en = 1'd0;
        pd80_clk = 1'd0;
        pd80_reset = 1'd0;
        pd81_in = 1'd0;
        pd81_write_en = 1'd0;
        pd81_clk = 1'd0;
        pd81_reset = 1'd0;
        pd82_in = 1'd0;
        pd82_write_en = 1'd0;
        pd82_clk = 1'd0;
        pd82_reset = 1'd0;
        pd83_in = 1'd0;
        pd83_write_en = 1'd0;
        pd83_clk = 1'd0;
        pd83_reset = 1'd0;
        pd84_in = 1'd0;
        pd84_write_en = 1'd0;
        pd84_clk = 1'd0;
        pd84_reset = 1'd0;
        pd85_in = 1'd0;
        pd85_write_en = 1'd0;
        pd85_clk = 1'd0;
        pd85_reset = 1'd0;
        pd86_in = 1'd0;
        pd86_write_en = 1'd0;
        pd86_clk = 1'd0;
        pd86_reset = 1'd0;
        pd87_in = 1'd0;
        pd87_write_en = 1'd0;
        pd87_clk = 1'd0;
        pd87_reset = 1'd0;
        pd88_in = 1'd0;
        pd88_write_en = 1'd0;
        pd88_clk = 1'd0;
        pd88_reset = 1'd0;
        pd89_in = 1'd0;
        pd89_write_en = 1'd0;
        pd89_clk = 1'd0;
        pd89_reset = 1'd0;
        pd90_in = 1'd0;
        pd90_write_en = 1'd0;
        pd90_clk = 1'd0;
        pd90_reset = 1'd0;
        pd91_in = 1'd0;
        pd91_write_en = 1'd0;
        pd91_clk = 1'd0;
        pd91_reset = 1'd0;
        pd92_in = 1'd0;
        pd92_write_en = 1'd0;
        pd92_clk = 1'd0;
        pd92_reset = 1'd0;
        fsm31_in = 3'd0;
        fsm31_write_en = 1'd0;
        fsm31_clk = 1'd0;
        fsm31_reset = 1'd0;
        pd93_in = 1'd0;
        pd93_write_en = 1'd0;
        pd93_clk = 1'd0;
        pd93_reset = 1'd0;
        fsm32_in = 4'd0;
        fsm32_write_en = 1'd0;
        fsm32_clk = 1'd0;
        fsm32_reset = 1'd0;
        pd94_in = 1'd0;
        pd94_write_en = 1'd0;
        pd94_clk = 1'd0;
        pd94_reset = 1'd0;
        fsm33_in = 1'd0;
        fsm33_write_en = 1'd0;
        fsm33_clk = 1'd0;
        fsm33_reset = 1'd0;
        write_zero_go_in = 1'd0;
        write_zero_done_in = 1'd0;
        write0_go_in = 1'd0;
        write0_done_in = 1'd0;
        write1_go_in = 1'd0;
        write1_done_in = 1'd0;
        write2_go_in = 1'd0;
        write2_done_in = 1'd0;
        write3_go_in = 1'd0;
        write3_done_in = 1'd0;
        write4_go_in = 1'd0;
        write4_done_in = 1'd0;
        write5_go_in = 1'd0;
        write5_done_in = 1'd0;
        write6_go_in = 1'd0;
        write6_done_in = 1'd0;
        write7_go_in = 1'd0;
        write7_done_in = 1'd0;
        write8_go_in = 1'd0;
        write8_done_in = 1'd0;
        write9_go_in = 1'd0;
        write9_done_in = 1'd0;
        write10_go_in = 1'd0;
        write10_done_in = 1'd0;
        write11_go_in = 1'd0;
        write11_done_in = 1'd0;
        write12_go_in = 1'd0;
        write12_done_in = 1'd0;
        write13_go_in = 1'd0;
        write13_done_in = 1'd0;
        write14_go_in = 1'd0;
        write14_done_in = 1'd0;
        write15_go_in = 1'd0;
        write15_done_in = 1'd0;
        write16_go_in = 1'd0;
        write16_done_in = 1'd0;
        write17_go_in = 1'd0;
        write17_done_in = 1'd0;
        write18_go_in = 1'd0;
        write18_done_in = 1'd0;
        write19_go_in = 1'd0;
        write19_done_in = 1'd0;
        write20_go_in = 1'd0;
        write20_done_in = 1'd0;
        write21_go_in = 1'd0;
        write21_done_in = 1'd0;
        write22_go_in = 1'd0;
        write22_done_in = 1'd0;
        write23_go_in = 1'd0;
        write23_done_in = 1'd0;
        write24_go_in = 1'd0;
        write24_done_in = 1'd0;
        write25_go_in = 1'd0;
        write25_done_in = 1'd0;
        write26_go_in = 1'd0;
        write26_done_in = 1'd0;
        write27_go_in = 1'd0;
        write27_done_in = 1'd0;
        write28_go_in = 1'd0;
        write28_done_in = 1'd0;
        write29_go_in = 1'd0;
        write29_done_in = 1'd0;
        write30_go_in = 1'd0;
        write30_done_in = 1'd0;
        write31_go_in = 1'd0;
        write31_done_in = 1'd0;
        find_write_index_go_in = 1'd0;
        find_write_index_done_in = 1'd0;
        default_to_zero_length_index_go_in = 1'd0;
        default_to_zero_length_index_done_in = 1'd0;
        save_index_go_in = 1'd0;
        save_index_done_in = 1'd0;
        is_length_zero0_go_in = 1'd0;
        is_length_zero0_done_in = 1'd0;
        invoke_go_in = 1'd0;
        invoke_done_in = 1'd0;
        invoke0_go_in = 1'd0;
        invoke0_done_in = 1'd0;
        invoke1_go_in = 1'd0;
        invoke1_done_in = 1'd0;
        invoke2_go_in = 1'd0;
        invoke2_done_in = 1'd0;
        invoke3_go_in = 1'd0;
        invoke3_done_in = 1'd0;
        invoke4_go_in = 1'd0;
        invoke4_done_in = 1'd0;
        invoke5_go_in = 1'd0;
        invoke5_done_in = 1'd0;
        invoke6_go_in = 1'd0;
        invoke6_done_in = 1'd0;
        invoke7_go_in = 1'd0;
        invoke7_done_in = 1'd0;
        invoke8_go_in = 1'd0;
        invoke8_done_in = 1'd0;
        invoke9_go_in = 1'd0;
        invoke9_done_in = 1'd0;
        invoke10_go_in = 1'd0;
        invoke10_done_in = 1'd0;
        invoke11_go_in = 1'd0;
        invoke11_done_in = 1'd0;
        invoke12_go_in = 1'd0;
        invoke12_done_in = 1'd0;
        invoke13_go_in = 1'd0;
        invoke13_done_in = 1'd0;
        invoke14_go_in = 1'd0;
        invoke14_done_in = 1'd0;
        invoke15_go_in = 1'd0;
        invoke15_done_in = 1'd0;
        invoke16_go_in = 1'd0;
        invoke16_done_in = 1'd0;
        invoke17_go_in = 1'd0;
        invoke17_done_in = 1'd0;
        invoke18_go_in = 1'd0;
        invoke18_done_in = 1'd0;
        invoke19_go_in = 1'd0;
        invoke19_done_in = 1'd0;
        invoke20_go_in = 1'd0;
        invoke20_done_in = 1'd0;
        invoke21_go_in = 1'd0;
        invoke21_done_in = 1'd0;
        invoke22_go_in = 1'd0;
        invoke22_done_in = 1'd0;
        invoke23_go_in = 1'd0;
        invoke23_done_in = 1'd0;
        invoke24_go_in = 1'd0;
        invoke24_done_in = 1'd0;
        invoke25_go_in = 1'd0;
        invoke25_done_in = 1'd0;
        invoke26_go_in = 1'd0;
        invoke26_done_in = 1'd0;
        invoke27_go_in = 1'd0;
        invoke27_done_in = 1'd0;
        invoke28_go_in = 1'd0;
        invoke28_done_in = 1'd0;
        invoke29_go_in = 1'd0;
        invoke29_done_in = 1'd0;
        invoke30_go_in = 1'd0;
        invoke30_done_in = 1'd0;
        invoke31_go_in = 1'd0;
        invoke31_done_in = 1'd0;
        invoke32_go_in = 1'd0;
        invoke32_done_in = 1'd0;
        invoke33_go_in = 1'd0;
        invoke33_done_in = 1'd0;
        invoke34_go_in = 1'd0;
        invoke34_done_in = 1'd0;
        invoke35_go_in = 1'd0;
        invoke35_done_in = 1'd0;
        invoke36_go_in = 1'd0;
        invoke36_done_in = 1'd0;
        invoke37_go_in = 1'd0;
        invoke37_done_in = 1'd0;
        invoke38_go_in = 1'd0;
        invoke38_done_in = 1'd0;
        invoke39_go_in = 1'd0;
        invoke39_done_in = 1'd0;
        invoke40_go_in = 1'd0;
        invoke40_done_in = 1'd0;
        invoke41_go_in = 1'd0;
        invoke41_done_in = 1'd0;
        invoke42_go_in = 1'd0;
        invoke42_done_in = 1'd0;
        invoke43_go_in = 1'd0;
        invoke43_done_in = 1'd0;
        invoke44_go_in = 1'd0;
        invoke44_done_in = 1'd0;
        invoke45_go_in = 1'd0;
        invoke45_done_in = 1'd0;
        invoke46_go_in = 1'd0;
        invoke46_done_in = 1'd0;
        invoke47_go_in = 1'd0;
        invoke47_done_in = 1'd0;
        invoke48_go_in = 1'd0;
        invoke48_done_in = 1'd0;
        invoke49_go_in = 1'd0;
        invoke49_done_in = 1'd0;
        invoke50_go_in = 1'd0;
        invoke50_done_in = 1'd0;
        invoke51_go_in = 1'd0;
        invoke51_done_in = 1'd0;
        invoke52_go_in = 1'd0;
        invoke52_done_in = 1'd0;
        invoke53_go_in = 1'd0;
        invoke53_done_in = 1'd0;
        invoke54_go_in = 1'd0;
        invoke54_done_in = 1'd0;
        invoke55_go_in = 1'd0;
        invoke55_done_in = 1'd0;
        invoke56_go_in = 1'd0;
        invoke56_done_in = 1'd0;
        invoke57_go_in = 1'd0;
        invoke57_done_in = 1'd0;
        invoke58_go_in = 1'd0;
        invoke58_done_in = 1'd0;
        invoke59_go_in = 1'd0;
        invoke59_done_in = 1'd0;
        invoke60_go_in = 1'd0;
        invoke60_done_in = 1'd0;
        invoke61_go_in = 1'd0;
        invoke61_done_in = 1'd0;
        par_go_in = 1'd0;
        par_done_in = 1'd0;
        tdcc_go_in = 1'd0;
        tdcc_done_in = 1'd0;
        tdcc0_go_in = 1'd0;
        tdcc0_done_in = 1'd0;
        tdcc1_go_in = 1'd0;
        tdcc1_done_in = 1'd0;
        tdcc2_go_in = 1'd0;
        tdcc2_done_in = 1'd0;
        tdcc3_go_in = 1'd0;
        tdcc3_done_in = 1'd0;
        tdcc4_go_in = 1'd0;
        tdcc4_done_in = 1'd0;
        tdcc5_go_in = 1'd0;
        tdcc5_done_in = 1'd0;
        tdcc6_go_in = 1'd0;
        tdcc6_done_in = 1'd0;
        tdcc7_go_in = 1'd0;
        tdcc7_done_in = 1'd0;
        tdcc8_go_in = 1'd0;
        tdcc8_done_in = 1'd0;
        tdcc9_go_in = 1'd0;
        tdcc9_done_in = 1'd0;
        tdcc10_go_in = 1'd0;
        tdcc10_done_in = 1'd0;
        tdcc11_go_in = 1'd0;
        tdcc11_done_in = 1'd0;
        tdcc12_go_in = 1'd0;
        tdcc12_done_in = 1'd0;
        tdcc13_go_in = 1'd0;
        tdcc13_done_in = 1'd0;
        tdcc14_go_in = 1'd0;
        tdcc14_done_in = 1'd0;
        tdcc15_go_in = 1'd0;
        tdcc15_done_in = 1'd0;
        tdcc16_go_in = 1'd0;
        tdcc16_done_in = 1'd0;
        tdcc17_go_in = 1'd0;
        tdcc17_done_in = 1'd0;
        tdcc18_go_in = 1'd0;
        tdcc18_done_in = 1'd0;
        tdcc19_go_in = 1'd0;
        tdcc19_done_in = 1'd0;
        tdcc20_go_in = 1'd0;
        tdcc20_done_in = 1'd0;
        tdcc21_go_in = 1'd0;
        tdcc21_done_in = 1'd0;
        tdcc22_go_in = 1'd0;
        tdcc22_done_in = 1'd0;
        tdcc23_go_in = 1'd0;
        tdcc23_done_in = 1'd0;
        tdcc24_go_in = 1'd0;
        tdcc24_done_in = 1'd0;
        tdcc25_go_in = 1'd0;
        tdcc25_done_in = 1'd0;
        tdcc26_go_in = 1'd0;
        tdcc26_done_in = 1'd0;
        tdcc27_go_in = 1'd0;
        tdcc27_done_in = 1'd0;
        tdcc28_go_in = 1'd0;
        tdcc28_done_in = 1'd0;
        tdcc29_go_in = 1'd0;
        tdcc29_done_in = 1'd0;
        tdcc30_go_in = 1'd0;
        tdcc30_done_in = 1'd0;
        par0_go_in = 1'd0;
        par0_done_in = 1'd0;
        par1_go_in = 1'd0;
        par1_done_in = 1'd0;
        par2_go_in = 1'd0;
        par2_done_in = 1'd0;
        par3_go_in = 1'd0;
        par3_done_in = 1'd0;
        par4_go_in = 1'd0;
        par4_done_in = 1'd0;
        par5_go_in = 1'd0;
        par5_done_in = 1'd0;
        tdcc31_go_in = 1'd0;
        tdcc31_done_in = 1'd0;
        tdcc32_go_in = 1'd0;
        tdcc32_done_in = 1'd0;
        tdcc33_go_in = 1'd0;
        tdcc33_done_in = 1'd0;
    end
    std_reg # (
        .WIDTH(32)
    ) p0 (
        .clk(p0_clk),
        .done(p0_done),
        .in(p0_in),
        .out(p0_out),
        .reset(p0_reset),
        .write_en(p0_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p1 (
        .clk(p1_clk),
        .done(p1_done),
        .in(p1_in),
        .out(p1_out),
        .reset(p1_reset),
        .write_en(p1_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p2 (
        .clk(p2_clk),
        .done(p2_done),
        .in(p2_in),
        .out(p2_out),
        .reset(p2_reset),
        .write_en(p2_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p3 (
        .clk(p3_clk),
        .done(p3_done),
        .in(p3_in),
        .out(p3_out),
        .reset(p3_reset),
        .write_en(p3_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p4 (
        .clk(p4_clk),
        .done(p4_done),
        .in(p4_in),
        .out(p4_out),
        .reset(p4_reset),
        .write_en(p4_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p5 (
        .clk(p5_clk),
        .done(p5_done),
        .in(p5_in),
        .out(p5_out),
        .reset(p5_reset),
        .write_en(p5_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p6 (
        .clk(p6_clk),
        .done(p6_done),
        .in(p6_in),
        .out(p6_out),
        .reset(p6_reset),
        .write_en(p6_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p7 (
        .clk(p7_clk),
        .done(p7_done),
        .in(p7_in),
        .out(p7_out),
        .reset(p7_reset),
        .write_en(p7_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p8 (
        .clk(p8_clk),
        .done(p8_done),
        .in(p8_in),
        .out(p8_out),
        .reset(p8_reset),
        .write_en(p8_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p9 (
        .clk(p9_clk),
        .done(p9_done),
        .in(p9_in),
        .out(p9_out),
        .reset(p9_reset),
        .write_en(p9_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p10 (
        .clk(p10_clk),
        .done(p10_done),
        .in(p10_in),
        .out(p10_out),
        .reset(p10_reset),
        .write_en(p10_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p11 (
        .clk(p11_clk),
        .done(p11_done),
        .in(p11_in),
        .out(p11_out),
        .reset(p11_reset),
        .write_en(p11_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p12 (
        .clk(p12_clk),
        .done(p12_done),
        .in(p12_in),
        .out(p12_out),
        .reset(p12_reset),
        .write_en(p12_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p13 (
        .clk(p13_clk),
        .done(p13_done),
        .in(p13_in),
        .out(p13_out),
        .reset(p13_reset),
        .write_en(p13_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p14 (
        .clk(p14_clk),
        .done(p14_done),
        .in(p14_in),
        .out(p14_out),
        .reset(p14_reset),
        .write_en(p14_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p15 (
        .clk(p15_clk),
        .done(p15_done),
        .in(p15_in),
        .out(p15_out),
        .reset(p15_reset),
        .write_en(p15_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p16 (
        .clk(p16_clk),
        .done(p16_done),
        .in(p16_in),
        .out(p16_out),
        .reset(p16_reset),
        .write_en(p16_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p17 (
        .clk(p17_clk),
        .done(p17_done),
        .in(p17_in),
        .out(p17_out),
        .reset(p17_reset),
        .write_en(p17_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p18 (
        .clk(p18_clk),
        .done(p18_done),
        .in(p18_in),
        .out(p18_out),
        .reset(p18_reset),
        .write_en(p18_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p19 (
        .clk(p19_clk),
        .done(p19_done),
        .in(p19_in),
        .out(p19_out),
        .reset(p19_reset),
        .write_en(p19_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p20 (
        .clk(p20_clk),
        .done(p20_done),
        .in(p20_in),
        .out(p20_out),
        .reset(p20_reset),
        .write_en(p20_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p21 (
        .clk(p21_clk),
        .done(p21_done),
        .in(p21_in),
        .out(p21_out),
        .reset(p21_reset),
        .write_en(p21_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p22 (
        .clk(p22_clk),
        .done(p22_done),
        .in(p22_in),
        .out(p22_out),
        .reset(p22_reset),
        .write_en(p22_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p23 (
        .clk(p23_clk),
        .done(p23_done),
        .in(p23_in),
        .out(p23_out),
        .reset(p23_reset),
        .write_en(p23_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p24 (
        .clk(p24_clk),
        .done(p24_done),
        .in(p24_in),
        .out(p24_out),
        .reset(p24_reset),
        .write_en(p24_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p25 (
        .clk(p25_clk),
        .done(p25_done),
        .in(p25_in),
        .out(p25_out),
        .reset(p25_reset),
        .write_en(p25_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p26 (
        .clk(p26_clk),
        .done(p26_done),
        .in(p26_in),
        .out(p26_out),
        .reset(p26_reset),
        .write_en(p26_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p27 (
        .clk(p27_clk),
        .done(p27_done),
        .in(p27_in),
        .out(p27_out),
        .reset(p27_reset),
        .write_en(p27_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p28 (
        .clk(p28_clk),
        .done(p28_done),
        .in(p28_in),
        .out(p28_out),
        .reset(p28_reset),
        .write_en(p28_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p29 (
        .clk(p29_clk),
        .done(p29_done),
        .in(p29_in),
        .out(p29_out),
        .reset(p29_reset),
        .write_en(p29_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p30 (
        .clk(p30_clk),
        .done(p30_done),
        .in(p30_in),
        .out(p30_out),
        .reset(p30_reset),
        .write_en(p30_write_en)
    );
    std_reg # (
        .WIDTH(32)
    ) p31 (
        .clk(p31_clk),
        .done(p31_done),
        .in(p31_in),
        .out(p31_out),
        .reset(p31_reset),
        .write_en(p31_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l0 (
        .clk(l0_clk),
        .done(l0_done),
        .in(l0_in),
        .out(l0_out),
        .reset(l0_reset),
        .write_en(l0_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l1 (
        .clk(l1_clk),
        .done(l1_done),
        .in(l1_in),
        .out(l1_out),
        .reset(l1_reset),
        .write_en(l1_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l2 (
        .clk(l2_clk),
        .done(l2_done),
        .in(l2_in),
        .out(l2_out),
        .reset(l2_reset),
        .write_en(l2_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l3 (
        .clk(l3_clk),
        .done(l3_done),
        .in(l3_in),
        .out(l3_out),
        .reset(l3_reset),
        .write_en(l3_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l4 (
        .clk(l4_clk),
        .done(l4_done),
        .in(l4_in),
        .out(l4_out),
        .reset(l4_reset),
        .write_en(l4_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l5 (
        .clk(l5_clk),
        .done(l5_done),
        .in(l5_in),
        .out(l5_out),
        .reset(l5_reset),
        .write_en(l5_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l6 (
        .clk(l6_clk),
        .done(l6_done),
        .in(l6_in),
        .out(l6_out),
        .reset(l6_reset),
        .write_en(l6_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l7 (
        .clk(l7_clk),
        .done(l7_done),
        .in(l7_in),
        .out(l7_out),
        .reset(l7_reset),
        .write_en(l7_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l8 (
        .clk(l8_clk),
        .done(l8_done),
        .in(l8_in),
        .out(l8_out),
        .reset(l8_reset),
        .write_en(l8_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l9 (
        .clk(l9_clk),
        .done(l9_done),
        .in(l9_in),
        .out(l9_out),
        .reset(l9_reset),
        .write_en(l9_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l10 (
        .clk(l10_clk),
        .done(l10_done),
        .in(l10_in),
        .out(l10_out),
        .reset(l10_reset),
        .write_en(l10_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l11 (
        .clk(l11_clk),
        .done(l11_done),
        .in(l11_in),
        .out(l11_out),
        .reset(l11_reset),
        .write_en(l11_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l12 (
        .clk(l12_clk),
        .done(l12_done),
        .in(l12_in),
        .out(l12_out),
        .reset(l12_reset),
        .write_en(l12_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l13 (
        .clk(l13_clk),
        .done(l13_done),
        .in(l13_in),
        .out(l13_out),
        .reset(l13_reset),
        .write_en(l13_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l14 (
        .clk(l14_clk),
        .done(l14_done),
        .in(l14_in),
        .out(l14_out),
        .reset(l14_reset),
        .write_en(l14_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l15 (
        .clk(l15_clk),
        .done(l15_done),
        .in(l15_in),
        .out(l15_out),
        .reset(l15_reset),
        .write_en(l15_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l16 (
        .clk(l16_clk),
        .done(l16_done),
        .in(l16_in),
        .out(l16_out),
        .reset(l16_reset),
        .write_en(l16_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l17 (
        .clk(l17_clk),
        .done(l17_done),
        .in(l17_in),
        .out(l17_out),
        .reset(l17_reset),
        .write_en(l17_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l18 (
        .clk(l18_clk),
        .done(l18_done),
        .in(l18_in),
        .out(l18_out),
        .reset(l18_reset),
        .write_en(l18_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l19 (
        .clk(l19_clk),
        .done(l19_done),
        .in(l19_in),
        .out(l19_out),
        .reset(l19_reset),
        .write_en(l19_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l20 (
        .clk(l20_clk),
        .done(l20_done),
        .in(l20_in),
        .out(l20_out),
        .reset(l20_reset),
        .write_en(l20_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l21 (
        .clk(l21_clk),
        .done(l21_done),
        .in(l21_in),
        .out(l21_out),
        .reset(l21_reset),
        .write_en(l21_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l22 (
        .clk(l22_clk),
        .done(l22_done),
        .in(l22_in),
        .out(l22_out),
        .reset(l22_reset),
        .write_en(l22_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l23 (
        .clk(l23_clk),
        .done(l23_done),
        .in(l23_in),
        .out(l23_out),
        .reset(l23_reset),
        .write_en(l23_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l24 (
        .clk(l24_clk),
        .done(l24_done),
        .in(l24_in),
        .out(l24_out),
        .reset(l24_reset),
        .write_en(l24_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l25 (
        .clk(l25_clk),
        .done(l25_done),
        .in(l25_in),
        .out(l25_out),
        .reset(l25_reset),
        .write_en(l25_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l26 (
        .clk(l26_clk),
        .done(l26_done),
        .in(l26_in),
        .out(l26_out),
        .reset(l26_reset),
        .write_en(l26_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l27 (
        .clk(l27_clk),
        .done(l27_done),
        .in(l27_in),
        .out(l27_out),
        .reset(l27_reset),
        .write_en(l27_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l28 (
        .clk(l28_clk),
        .done(l28_done),
        .in(l28_in),
        .out(l28_out),
        .reset(l28_reset),
        .write_en(l28_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l29 (
        .clk(l29_clk),
        .done(l29_done),
        .in(l29_in),
        .out(l29_out),
        .reset(l29_reset),
        .write_en(l29_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l30 (
        .clk(l30_clk),
        .done(l30_done),
        .in(l30_in),
        .out(l30_out),
        .reset(l30_reset),
        .write_en(l30_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) l31 (
        .clk(l31_clk),
        .done(l31_done),
        .in(l31_in),
        .out(l31_out),
        .reset(l31_reset),
        .write_en(l31_write_en)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index0 (
        .left(is_index0_left),
        .out(is_index0_out),
        .right(is_index0_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index1 (
        .left(is_index1_left),
        .out(is_index1_out),
        .right(is_index1_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index2 (
        .left(is_index2_left),
        .out(is_index2_out),
        .right(is_index2_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index3 (
        .left(is_index3_left),
        .out(is_index3_out),
        .right(is_index3_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index4 (
        .left(is_index4_left),
        .out(is_index4_out),
        .right(is_index4_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index5 (
        .left(is_index5_left),
        .out(is_index5_out),
        .right(is_index5_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index6 (
        .left(is_index6_left),
        .out(is_index6_out),
        .right(is_index6_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index7 (
        .left(is_index7_left),
        .out(is_index7_out),
        .right(is_index7_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index8 (
        .left(is_index8_left),
        .out(is_index8_out),
        .right(is_index8_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index9 (
        .left(is_index9_left),
        .out(is_index9_out),
        .right(is_index9_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index10 (
        .left(is_index10_left),
        .out(is_index10_out),
        .right(is_index10_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index11 (
        .left(is_index11_left),
        .out(is_index11_out),
        .right(is_index11_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index12 (
        .left(is_index12_left),
        .out(is_index12_out),
        .right(is_index12_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index13 (
        .left(is_index13_left),
        .out(is_index13_out),
        .right(is_index13_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index14 (
        .left(is_index14_left),
        .out(is_index14_out),
        .right(is_index14_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index15 (
        .left(is_index15_left),
        .out(is_index15_out),
        .right(is_index15_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index16 (
        .left(is_index16_left),
        .out(is_index16_out),
        .right(is_index16_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index17 (
        .left(is_index17_left),
        .out(is_index17_out),
        .right(is_index17_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index18 (
        .left(is_index18_left),
        .out(is_index18_out),
        .right(is_index18_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index19 (
        .left(is_index19_left),
        .out(is_index19_out),
        .right(is_index19_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index20 (
        .left(is_index20_left),
        .out(is_index20_out),
        .right(is_index20_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index21 (
        .left(is_index21_left),
        .out(is_index21_out),
        .right(is_index21_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index22 (
        .left(is_index22_left),
        .out(is_index22_out),
        .right(is_index22_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index23 (
        .left(is_index23_left),
        .out(is_index23_out),
        .right(is_index23_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index24 (
        .left(is_index24_left),
        .out(is_index24_out),
        .right(is_index24_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index25 (
        .left(is_index25_left),
        .out(is_index25_out),
        .right(is_index25_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index26 (
        .left(is_index26_left),
        .out(is_index26_out),
        .right(is_index26_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index27 (
        .left(is_index27_left),
        .out(is_index27_out),
        .right(is_index27_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index28 (
        .left(is_index28_left),
        .out(is_index28_out),
        .right(is_index28_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index29 (
        .left(is_index29_left),
        .out(is_index29_out),
        .right(is_index29_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index30 (
        .left(is_index30_left),
        .out(is_index30_out),
        .right(is_index30_right)
    );
    std_eq # (
        .WIDTH(5)
    ) is_index31 (
        .left(is_index31_left),
        .out(is_index31_out),
        .right(is_index31_right)
    );
    std_reg # (
        .WIDTH(5)
    ) zero_index (
        .clk(zero_index_clk),
        .done(zero_index_done),
        .in(zero_index_in),
        .out(zero_index_out),
        .reset(zero_index_reset),
        .write_en(zero_index_write_en)
    );
    std_eq # (
        .WIDTH(6)
    ) z_eq (
        .left(z_eq_left),
        .out(z_eq_out),
        .right(z_eq_right)
    );
    std_slice # (
        .IN_WIDTH(6),
        .OUT_WIDTH(5)
    ) slice (
        .in(slice_in),
        .out(slice_out)
    );
    std_sub # (
        .WIDTH(6)
    ) sub (
        .left(sub_left),
        .out(sub_out),
        .right(sub_right)
    );
    match_element me0 (
        .clk(me0_clk),
        .done(me0_done),
        .go(me0_go),
        .in(me0_in),
        .length(me0_length),
        .out(me0_out),
        .prefix(me0_prefix),
        .reset(me0_reset)
    );
    match_element me1 (
        .clk(me1_clk),
        .done(me1_done),
        .go(me1_go),
        .in(me1_in),
        .length(me1_length),
        .out(me1_out),
        .prefix(me1_prefix),
        .reset(me1_reset)
    );
    match_element me2 (
        .clk(me2_clk),
        .done(me2_done),
        .go(me2_go),
        .in(me2_in),
        .length(me2_length),
        .out(me2_out),
        .prefix(me2_prefix),
        .reset(me2_reset)
    );
    match_element me3 (
        .clk(me3_clk),
        .done(me3_done),
        .go(me3_go),
        .in(me3_in),
        .length(me3_length),
        .out(me3_out),
        .prefix(me3_prefix),
        .reset(me3_reset)
    );
    match_element me4 (
        .clk(me4_clk),
        .done(me4_done),
        .go(me4_go),
        .in(me4_in),
        .length(me4_length),
        .out(me4_out),
        .prefix(me4_prefix),
        .reset(me4_reset)
    );
    match_element me5 (
        .clk(me5_clk),
        .done(me5_done),
        .go(me5_go),
        .in(me5_in),
        .length(me5_length),
        .out(me5_out),
        .prefix(me5_prefix),
        .reset(me5_reset)
    );
    match_element me6 (
        .clk(me6_clk),
        .done(me6_done),
        .go(me6_go),
        .in(me6_in),
        .length(me6_length),
        .out(me6_out),
        .prefix(me6_prefix),
        .reset(me6_reset)
    );
    match_element me7 (
        .clk(me7_clk),
        .done(me7_done),
        .go(me7_go),
        .in(me7_in),
        .length(me7_length),
        .out(me7_out),
        .prefix(me7_prefix),
        .reset(me7_reset)
    );
    match_element me8 (
        .clk(me8_clk),
        .done(me8_done),
        .go(me8_go),
        .in(me8_in),
        .length(me8_length),
        .out(me8_out),
        .prefix(me8_prefix),
        .reset(me8_reset)
    );
    match_element me9 (
        .clk(me9_clk),
        .done(me9_done),
        .go(me9_go),
        .in(me9_in),
        .length(me9_length),
        .out(me9_out),
        .prefix(me9_prefix),
        .reset(me9_reset)
    );
    match_element me10 (
        .clk(me10_clk),
        .done(me10_done),
        .go(me10_go),
        .in(me10_in),
        .length(me10_length),
        .out(me10_out),
        .prefix(me10_prefix),
        .reset(me10_reset)
    );
    match_element me11 (
        .clk(me11_clk),
        .done(me11_done),
        .go(me11_go),
        .in(me11_in),
        .length(me11_length),
        .out(me11_out),
        .prefix(me11_prefix),
        .reset(me11_reset)
    );
    match_element me12 (
        .clk(me12_clk),
        .done(me12_done),
        .go(me12_go),
        .in(me12_in),
        .length(me12_length),
        .out(me12_out),
        .prefix(me12_prefix),
        .reset(me12_reset)
    );
    match_element me13 (
        .clk(me13_clk),
        .done(me13_done),
        .go(me13_go),
        .in(me13_in),
        .length(me13_length),
        .out(me13_out),
        .prefix(me13_prefix),
        .reset(me13_reset)
    );
    match_element me14 (
        .clk(me14_clk),
        .done(me14_done),
        .go(me14_go),
        .in(me14_in),
        .length(me14_length),
        .out(me14_out),
        .prefix(me14_prefix),
        .reset(me14_reset)
    );
    match_element me15 (
        .clk(me15_clk),
        .done(me15_done),
        .go(me15_go),
        .in(me15_in),
        .length(me15_length),
        .out(me15_out),
        .prefix(me15_prefix),
        .reset(me15_reset)
    );
    match_element me16 (
        .clk(me16_clk),
        .done(me16_done),
        .go(me16_go),
        .in(me16_in),
        .length(me16_length),
        .out(me16_out),
        .prefix(me16_prefix),
        .reset(me16_reset)
    );
    match_element me17 (
        .clk(me17_clk),
        .done(me17_done),
        .go(me17_go),
        .in(me17_in),
        .length(me17_length),
        .out(me17_out),
        .prefix(me17_prefix),
        .reset(me17_reset)
    );
    match_element me18 (
        .clk(me18_clk),
        .done(me18_done),
        .go(me18_go),
        .in(me18_in),
        .length(me18_length),
        .out(me18_out),
        .prefix(me18_prefix),
        .reset(me18_reset)
    );
    match_element me19 (
        .clk(me19_clk),
        .done(me19_done),
        .go(me19_go),
        .in(me19_in),
        .length(me19_length),
        .out(me19_out),
        .prefix(me19_prefix),
        .reset(me19_reset)
    );
    match_element me20 (
        .clk(me20_clk),
        .done(me20_done),
        .go(me20_go),
        .in(me20_in),
        .length(me20_length),
        .out(me20_out),
        .prefix(me20_prefix),
        .reset(me20_reset)
    );
    match_element me21 (
        .clk(me21_clk),
        .done(me21_done),
        .go(me21_go),
        .in(me21_in),
        .length(me21_length),
        .out(me21_out),
        .prefix(me21_prefix),
        .reset(me21_reset)
    );
    match_element me22 (
        .clk(me22_clk),
        .done(me22_done),
        .go(me22_go),
        .in(me22_in),
        .length(me22_length),
        .out(me22_out),
        .prefix(me22_prefix),
        .reset(me22_reset)
    );
    match_element me23 (
        .clk(me23_clk),
        .done(me23_done),
        .go(me23_go),
        .in(me23_in),
        .length(me23_length),
        .out(me23_out),
        .prefix(me23_prefix),
        .reset(me23_reset)
    );
    match_element me24 (
        .clk(me24_clk),
        .done(me24_done),
        .go(me24_go),
        .in(me24_in),
        .length(me24_length),
        .out(me24_out),
        .prefix(me24_prefix),
        .reset(me24_reset)
    );
    match_element me25 (
        .clk(me25_clk),
        .done(me25_done),
        .go(me25_go),
        .in(me25_in),
        .length(me25_length),
        .out(me25_out),
        .prefix(me25_prefix),
        .reset(me25_reset)
    );
    match_element me26 (
        .clk(me26_clk),
        .done(me26_done),
        .go(me26_go),
        .in(me26_in),
        .length(me26_length),
        .out(me26_out),
        .prefix(me26_prefix),
        .reset(me26_reset)
    );
    match_element me27 (
        .clk(me27_clk),
        .done(me27_done),
        .go(me27_go),
        .in(me27_in),
        .length(me27_length),
        .out(me27_out),
        .prefix(me27_prefix),
        .reset(me27_reset)
    );
    match_element me28 (
        .clk(me28_clk),
        .done(me28_done),
        .go(me28_go),
        .in(me28_in),
        .length(me28_length),
        .out(me28_out),
        .prefix(me28_prefix),
        .reset(me28_reset)
    );
    match_element me29 (
        .clk(me29_clk),
        .done(me29_done),
        .go(me29_go),
        .in(me29_in),
        .length(me29_length),
        .out(me29_out),
        .prefix(me29_prefix),
        .reset(me29_reset)
    );
    match_element me30 (
        .clk(me30_clk),
        .done(me30_done),
        .go(me30_go),
        .in(me30_in),
        .length(me30_length),
        .out(me30_out),
        .prefix(me30_prefix),
        .reset(me30_reset)
    );
    match_element me31 (
        .clk(me31_clk),
        .done(me31_done),
        .go(me31_go),
        .in(me31_in),
        .length(me31_length),
        .out(me31_out),
        .prefix(me31_prefix),
        .reset(me31_reset)
    );
    comparator_element ce00 (
        .addrA(ce00_addrA),
        .addrB(ce00_addrB),
        .addrX(ce00_addrX),
        .clk(ce00_clk),
        .done(ce00_done),
        .go(ce00_go),
        .lenA(ce00_lenA),
        .lenB(ce00_lenB),
        .lenX(ce00_lenX),
        .mlA(ce00_mlA),
        .mlB(ce00_mlB),
        .mlX(ce00_mlX),
        .reset(ce00_reset)
    );
    comparator_element ce01 (
        .addrA(ce01_addrA),
        .addrB(ce01_addrB),
        .addrX(ce01_addrX),
        .clk(ce01_clk),
        .done(ce01_done),
        .go(ce01_go),
        .lenA(ce01_lenA),
        .lenB(ce01_lenB),
        .lenX(ce01_lenX),
        .mlA(ce01_mlA),
        .mlB(ce01_mlB),
        .mlX(ce01_mlX),
        .reset(ce01_reset)
    );
    comparator_element ce02 (
        .addrA(ce02_addrA),
        .addrB(ce02_addrB),
        .addrX(ce02_addrX),
        .clk(ce02_clk),
        .done(ce02_done),
        .go(ce02_go),
        .lenA(ce02_lenA),
        .lenB(ce02_lenB),
        .lenX(ce02_lenX),
        .mlA(ce02_mlA),
        .mlB(ce02_mlB),
        .mlX(ce02_mlX),
        .reset(ce02_reset)
    );
    comparator_element ce03 (
        .addrA(ce03_addrA),
        .addrB(ce03_addrB),
        .addrX(ce03_addrX),
        .clk(ce03_clk),
        .done(ce03_done),
        .go(ce03_go),
        .lenA(ce03_lenA),
        .lenB(ce03_lenB),
        .lenX(ce03_lenX),
        .mlA(ce03_mlA),
        .mlB(ce03_mlB),
        .mlX(ce03_mlX),
        .reset(ce03_reset)
    );
    comparator_element ce04 (
        .addrA(ce04_addrA),
        .addrB(ce04_addrB),
        .addrX(ce04_addrX),
        .clk(ce04_clk),
        .done(ce04_done),
        .go(ce04_go),
        .lenA(ce04_lenA),
        .lenB(ce04_lenB),
        .lenX(ce04_lenX),
        .mlA(ce04_mlA),
        .mlB(ce04_mlB),
        .mlX(ce04_mlX),
        .reset(ce04_reset)
    );
    comparator_element ce05 (
        .addrA(ce05_addrA),
        .addrB(ce05_addrB),
        .addrX(ce05_addrX),
        .clk(ce05_clk),
        .done(ce05_done),
        .go(ce05_go),
        .lenA(ce05_lenA),
        .lenB(ce05_lenB),
        .lenX(ce05_lenX),
        .mlA(ce05_mlA),
        .mlB(ce05_mlB),
        .mlX(ce05_mlX),
        .reset(ce05_reset)
    );
    comparator_element ce06 (
        .addrA(ce06_addrA),
        .addrB(ce06_addrB),
        .addrX(ce06_addrX),
        .clk(ce06_clk),
        .done(ce06_done),
        .go(ce06_go),
        .lenA(ce06_lenA),
        .lenB(ce06_lenB),
        .lenX(ce06_lenX),
        .mlA(ce06_mlA),
        .mlB(ce06_mlB),
        .mlX(ce06_mlX),
        .reset(ce06_reset)
    );
    comparator_element ce07 (
        .addrA(ce07_addrA),
        .addrB(ce07_addrB),
        .addrX(ce07_addrX),
        .clk(ce07_clk),
        .done(ce07_done),
        .go(ce07_go),
        .lenA(ce07_lenA),
        .lenB(ce07_lenB),
        .lenX(ce07_lenX),
        .mlA(ce07_mlA),
        .mlB(ce07_mlB),
        .mlX(ce07_mlX),
        .reset(ce07_reset)
    );
    comparator_element ce08 (
        .addrA(ce08_addrA),
        .addrB(ce08_addrB),
        .addrX(ce08_addrX),
        .clk(ce08_clk),
        .done(ce08_done),
        .go(ce08_go),
        .lenA(ce08_lenA),
        .lenB(ce08_lenB),
        .lenX(ce08_lenX),
        .mlA(ce08_mlA),
        .mlB(ce08_mlB),
        .mlX(ce08_mlX),
        .reset(ce08_reset)
    );
    comparator_element ce09 (
        .addrA(ce09_addrA),
        .addrB(ce09_addrB),
        .addrX(ce09_addrX),
        .clk(ce09_clk),
        .done(ce09_done),
        .go(ce09_go),
        .lenA(ce09_lenA),
        .lenB(ce09_lenB),
        .lenX(ce09_lenX),
        .mlA(ce09_mlA),
        .mlB(ce09_mlB),
        .mlX(ce09_mlX),
        .reset(ce09_reset)
    );
    comparator_element ce010 (
        .addrA(ce010_addrA),
        .addrB(ce010_addrB),
        .addrX(ce010_addrX),
        .clk(ce010_clk),
        .done(ce010_done),
        .go(ce010_go),
        .lenA(ce010_lenA),
        .lenB(ce010_lenB),
        .lenX(ce010_lenX),
        .mlA(ce010_mlA),
        .mlB(ce010_mlB),
        .mlX(ce010_mlX),
        .reset(ce010_reset)
    );
    comparator_element ce011 (
        .addrA(ce011_addrA),
        .addrB(ce011_addrB),
        .addrX(ce011_addrX),
        .clk(ce011_clk),
        .done(ce011_done),
        .go(ce011_go),
        .lenA(ce011_lenA),
        .lenB(ce011_lenB),
        .lenX(ce011_lenX),
        .mlA(ce011_mlA),
        .mlB(ce011_mlB),
        .mlX(ce011_mlX),
        .reset(ce011_reset)
    );
    comparator_element ce012 (
        .addrA(ce012_addrA),
        .addrB(ce012_addrB),
        .addrX(ce012_addrX),
        .clk(ce012_clk),
        .done(ce012_done),
        .go(ce012_go),
        .lenA(ce012_lenA),
        .lenB(ce012_lenB),
        .lenX(ce012_lenX),
        .mlA(ce012_mlA),
        .mlB(ce012_mlB),
        .mlX(ce012_mlX),
        .reset(ce012_reset)
    );
    comparator_element ce013 (
        .addrA(ce013_addrA),
        .addrB(ce013_addrB),
        .addrX(ce013_addrX),
        .clk(ce013_clk),
        .done(ce013_done),
        .go(ce013_go),
        .lenA(ce013_lenA),
        .lenB(ce013_lenB),
        .lenX(ce013_lenX),
        .mlA(ce013_mlA),
        .mlB(ce013_mlB),
        .mlX(ce013_mlX),
        .reset(ce013_reset)
    );
    comparator_element ce014 (
        .addrA(ce014_addrA),
        .addrB(ce014_addrB),
        .addrX(ce014_addrX),
        .clk(ce014_clk),
        .done(ce014_done),
        .go(ce014_go),
        .lenA(ce014_lenA),
        .lenB(ce014_lenB),
        .lenX(ce014_lenX),
        .mlA(ce014_mlA),
        .mlB(ce014_mlB),
        .mlX(ce014_mlX),
        .reset(ce014_reset)
    );
    comparator_element ce015 (
        .addrA(ce015_addrA),
        .addrB(ce015_addrB),
        .addrX(ce015_addrX),
        .clk(ce015_clk),
        .done(ce015_done),
        .go(ce015_go),
        .lenA(ce015_lenA),
        .lenB(ce015_lenB),
        .lenX(ce015_lenX),
        .mlA(ce015_mlA),
        .mlB(ce015_mlB),
        .mlX(ce015_mlX),
        .reset(ce015_reset)
    );
    comparator_element ce10 (
        .addrA(ce10_addrA),
        .addrB(ce10_addrB),
        .addrX(ce10_addrX),
        .clk(ce10_clk),
        .done(ce10_done),
        .go(ce10_go),
        .lenA(ce10_lenA),
        .lenB(ce10_lenB),
        .lenX(ce10_lenX),
        .mlA(ce10_mlA),
        .mlB(ce10_mlB),
        .mlX(ce10_mlX),
        .reset(ce10_reset)
    );
    comparator_element ce11 (
        .addrA(ce11_addrA),
        .addrB(ce11_addrB),
        .addrX(ce11_addrX),
        .clk(ce11_clk),
        .done(ce11_done),
        .go(ce11_go),
        .lenA(ce11_lenA),
        .lenB(ce11_lenB),
        .lenX(ce11_lenX),
        .mlA(ce11_mlA),
        .mlB(ce11_mlB),
        .mlX(ce11_mlX),
        .reset(ce11_reset)
    );
    comparator_element ce12 (
        .addrA(ce12_addrA),
        .addrB(ce12_addrB),
        .addrX(ce12_addrX),
        .clk(ce12_clk),
        .done(ce12_done),
        .go(ce12_go),
        .lenA(ce12_lenA),
        .lenB(ce12_lenB),
        .lenX(ce12_lenX),
        .mlA(ce12_mlA),
        .mlB(ce12_mlB),
        .mlX(ce12_mlX),
        .reset(ce12_reset)
    );
    comparator_element ce13 (
        .addrA(ce13_addrA),
        .addrB(ce13_addrB),
        .addrX(ce13_addrX),
        .clk(ce13_clk),
        .done(ce13_done),
        .go(ce13_go),
        .lenA(ce13_lenA),
        .lenB(ce13_lenB),
        .lenX(ce13_lenX),
        .mlA(ce13_mlA),
        .mlB(ce13_mlB),
        .mlX(ce13_mlX),
        .reset(ce13_reset)
    );
    comparator_element ce14 (
        .addrA(ce14_addrA),
        .addrB(ce14_addrB),
        .addrX(ce14_addrX),
        .clk(ce14_clk),
        .done(ce14_done),
        .go(ce14_go),
        .lenA(ce14_lenA),
        .lenB(ce14_lenB),
        .lenX(ce14_lenX),
        .mlA(ce14_mlA),
        .mlB(ce14_mlB),
        .mlX(ce14_mlX),
        .reset(ce14_reset)
    );
    comparator_element ce15 (
        .addrA(ce15_addrA),
        .addrB(ce15_addrB),
        .addrX(ce15_addrX),
        .clk(ce15_clk),
        .done(ce15_done),
        .go(ce15_go),
        .lenA(ce15_lenA),
        .lenB(ce15_lenB),
        .lenX(ce15_lenX),
        .mlA(ce15_mlA),
        .mlB(ce15_mlB),
        .mlX(ce15_mlX),
        .reset(ce15_reset)
    );
    comparator_element ce16 (
        .addrA(ce16_addrA),
        .addrB(ce16_addrB),
        .addrX(ce16_addrX),
        .clk(ce16_clk),
        .done(ce16_done),
        .go(ce16_go),
        .lenA(ce16_lenA),
        .lenB(ce16_lenB),
        .lenX(ce16_lenX),
        .mlA(ce16_mlA),
        .mlB(ce16_mlB),
        .mlX(ce16_mlX),
        .reset(ce16_reset)
    );
    comparator_element ce17 (
        .addrA(ce17_addrA),
        .addrB(ce17_addrB),
        .addrX(ce17_addrX),
        .clk(ce17_clk),
        .done(ce17_done),
        .go(ce17_go),
        .lenA(ce17_lenA),
        .lenB(ce17_lenB),
        .lenX(ce17_lenX),
        .mlA(ce17_mlA),
        .mlB(ce17_mlB),
        .mlX(ce17_mlX),
        .reset(ce17_reset)
    );
    comparator_element ce20 (
        .addrA(ce20_addrA),
        .addrB(ce20_addrB),
        .addrX(ce20_addrX),
        .clk(ce20_clk),
        .done(ce20_done),
        .go(ce20_go),
        .lenA(ce20_lenA),
        .lenB(ce20_lenB),
        .lenX(ce20_lenX),
        .mlA(ce20_mlA),
        .mlB(ce20_mlB),
        .mlX(ce20_mlX),
        .reset(ce20_reset)
    );
    comparator_element ce21 (
        .addrA(ce21_addrA),
        .addrB(ce21_addrB),
        .addrX(ce21_addrX),
        .clk(ce21_clk),
        .done(ce21_done),
        .go(ce21_go),
        .lenA(ce21_lenA),
        .lenB(ce21_lenB),
        .lenX(ce21_lenX),
        .mlA(ce21_mlA),
        .mlB(ce21_mlB),
        .mlX(ce21_mlX),
        .reset(ce21_reset)
    );
    comparator_element ce22 (
        .addrA(ce22_addrA),
        .addrB(ce22_addrB),
        .addrX(ce22_addrX),
        .clk(ce22_clk),
        .done(ce22_done),
        .go(ce22_go),
        .lenA(ce22_lenA),
        .lenB(ce22_lenB),
        .lenX(ce22_lenX),
        .mlA(ce22_mlA),
        .mlB(ce22_mlB),
        .mlX(ce22_mlX),
        .reset(ce22_reset)
    );
    comparator_element ce23 (
        .addrA(ce23_addrA),
        .addrB(ce23_addrB),
        .addrX(ce23_addrX),
        .clk(ce23_clk),
        .done(ce23_done),
        .go(ce23_go),
        .lenA(ce23_lenA),
        .lenB(ce23_lenB),
        .lenX(ce23_lenX),
        .mlA(ce23_mlA),
        .mlB(ce23_mlB),
        .mlX(ce23_mlX),
        .reset(ce23_reset)
    );
    comparator_element ce30 (
        .addrA(ce30_addrA),
        .addrB(ce30_addrB),
        .addrX(ce30_addrX),
        .clk(ce30_clk),
        .done(ce30_done),
        .go(ce30_go),
        .lenA(ce30_lenA),
        .lenB(ce30_lenB),
        .lenX(ce30_lenX),
        .mlA(ce30_mlA),
        .mlB(ce30_mlB),
        .mlX(ce30_mlX),
        .reset(ce30_reset)
    );
    comparator_element ce31 (
        .addrA(ce31_addrA),
        .addrB(ce31_addrB),
        .addrX(ce31_addrX),
        .clk(ce31_clk),
        .done(ce31_done),
        .go(ce31_go),
        .lenA(ce31_lenA),
        .lenB(ce31_lenB),
        .lenX(ce31_lenX),
        .mlA(ce31_mlA),
        .mlB(ce31_mlB),
        .mlX(ce31_mlX),
        .reset(ce31_reset)
    );
    comparator_element ce40 (
        .addrA(ce40_addrA),
        .addrB(ce40_addrB),
        .addrX(ce40_addrX),
        .clk(ce40_clk),
        .done(ce40_done),
        .go(ce40_go),
        .lenA(ce40_lenA),
        .lenB(ce40_lenB),
        .lenX(ce40_lenX),
        .mlA(ce40_mlA),
        .mlB(ce40_mlB),
        .mlX(ce40_mlX),
        .reset(ce40_reset)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg0 (
        .clk(comb_reg0_clk),
        .done(comb_reg0_done),
        .in(comb_reg0_in),
        .out(comb_reg0_out),
        .reset(comb_reg0_reset),
        .write_en(comb_reg0_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg1 (
        .clk(comb_reg1_clk),
        .done(comb_reg1_done),
        .in(comb_reg1_in),
        .out(comb_reg1_out),
        .reset(comb_reg1_reset),
        .write_en(comb_reg1_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg2 (
        .clk(comb_reg2_clk),
        .done(comb_reg2_done),
        .in(comb_reg2_in),
        .out(comb_reg2_out),
        .reset(comb_reg2_reset),
        .write_en(comb_reg2_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg3 (
        .clk(comb_reg3_clk),
        .done(comb_reg3_done),
        .in(comb_reg3_in),
        .out(comb_reg3_out),
        .reset(comb_reg3_reset),
        .write_en(comb_reg3_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg4 (
        .clk(comb_reg4_clk),
        .done(comb_reg4_done),
        .in(comb_reg4_in),
        .out(comb_reg4_out),
        .reset(comb_reg4_reset),
        .write_en(comb_reg4_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg5 (
        .clk(comb_reg5_clk),
        .done(comb_reg5_done),
        .in(comb_reg5_in),
        .out(comb_reg5_out),
        .reset(comb_reg5_reset),
        .write_en(comb_reg5_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg6 (
        .clk(comb_reg6_clk),
        .done(comb_reg6_done),
        .in(comb_reg6_in),
        .out(comb_reg6_out),
        .reset(comb_reg6_reset),
        .write_en(comb_reg6_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg7 (
        .clk(comb_reg7_clk),
        .done(comb_reg7_done),
        .in(comb_reg7_in),
        .out(comb_reg7_out),
        .reset(comb_reg7_reset),
        .write_en(comb_reg7_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg8 (
        .clk(comb_reg8_clk),
        .done(comb_reg8_done),
        .in(comb_reg8_in),
        .out(comb_reg8_out),
        .reset(comb_reg8_reset),
        .write_en(comb_reg8_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg9 (
        .clk(comb_reg9_clk),
        .done(comb_reg9_done),
        .in(comb_reg9_in),
        .out(comb_reg9_out),
        .reset(comb_reg9_reset),
        .write_en(comb_reg9_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg10 (
        .clk(comb_reg10_clk),
        .done(comb_reg10_done),
        .in(comb_reg10_in),
        .out(comb_reg10_out),
        .reset(comb_reg10_reset),
        .write_en(comb_reg10_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg11 (
        .clk(comb_reg11_clk),
        .done(comb_reg11_done),
        .in(comb_reg11_in),
        .out(comb_reg11_out),
        .reset(comb_reg11_reset),
        .write_en(comb_reg11_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg12 (
        .clk(comb_reg12_clk),
        .done(comb_reg12_done),
        .in(comb_reg12_in),
        .out(comb_reg12_out),
        .reset(comb_reg12_reset),
        .write_en(comb_reg12_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg13 (
        .clk(comb_reg13_clk),
        .done(comb_reg13_done),
        .in(comb_reg13_in),
        .out(comb_reg13_out),
        .reset(comb_reg13_reset),
        .write_en(comb_reg13_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg14 (
        .clk(comb_reg14_clk),
        .done(comb_reg14_done),
        .in(comb_reg14_in),
        .out(comb_reg14_out),
        .reset(comb_reg14_reset),
        .write_en(comb_reg14_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg15 (
        .clk(comb_reg15_clk),
        .done(comb_reg15_done),
        .in(comb_reg15_in),
        .out(comb_reg15_out),
        .reset(comb_reg15_reset),
        .write_en(comb_reg15_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg16 (
        .clk(comb_reg16_clk),
        .done(comb_reg16_done),
        .in(comb_reg16_in),
        .out(comb_reg16_out),
        .reset(comb_reg16_reset),
        .write_en(comb_reg16_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg17 (
        .clk(comb_reg17_clk),
        .done(comb_reg17_done),
        .in(comb_reg17_in),
        .out(comb_reg17_out),
        .reset(comb_reg17_reset),
        .write_en(comb_reg17_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg18 (
        .clk(comb_reg18_clk),
        .done(comb_reg18_done),
        .in(comb_reg18_in),
        .out(comb_reg18_out),
        .reset(comb_reg18_reset),
        .write_en(comb_reg18_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg19 (
        .clk(comb_reg19_clk),
        .done(comb_reg19_done),
        .in(comb_reg19_in),
        .out(comb_reg19_out),
        .reset(comb_reg19_reset),
        .write_en(comb_reg19_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg20 (
        .clk(comb_reg20_clk),
        .done(comb_reg20_done),
        .in(comb_reg20_in),
        .out(comb_reg20_out),
        .reset(comb_reg20_reset),
        .write_en(comb_reg20_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg21 (
        .clk(comb_reg21_clk),
        .done(comb_reg21_done),
        .in(comb_reg21_in),
        .out(comb_reg21_out),
        .reset(comb_reg21_reset),
        .write_en(comb_reg21_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg22 (
        .clk(comb_reg22_clk),
        .done(comb_reg22_done),
        .in(comb_reg22_in),
        .out(comb_reg22_out),
        .reset(comb_reg22_reset),
        .write_en(comb_reg22_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg23 (
        .clk(comb_reg23_clk),
        .done(comb_reg23_done),
        .in(comb_reg23_in),
        .out(comb_reg23_out),
        .reset(comb_reg23_reset),
        .write_en(comb_reg23_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg24 (
        .clk(comb_reg24_clk),
        .done(comb_reg24_done),
        .in(comb_reg24_in),
        .out(comb_reg24_out),
        .reset(comb_reg24_reset),
        .write_en(comb_reg24_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg25 (
        .clk(comb_reg25_clk),
        .done(comb_reg25_done),
        .in(comb_reg25_in),
        .out(comb_reg25_out),
        .reset(comb_reg25_reset),
        .write_en(comb_reg25_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg26 (
        .clk(comb_reg26_clk),
        .done(comb_reg26_done),
        .in(comb_reg26_in),
        .out(comb_reg26_out),
        .reset(comb_reg26_reset),
        .write_en(comb_reg26_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg27 (
        .clk(comb_reg27_clk),
        .done(comb_reg27_done),
        .in(comb_reg27_in),
        .out(comb_reg27_out),
        .reset(comb_reg27_reset),
        .write_en(comb_reg27_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg28 (
        .clk(comb_reg28_clk),
        .done(comb_reg28_done),
        .in(comb_reg28_in),
        .out(comb_reg28_out),
        .reset(comb_reg28_reset),
        .write_en(comb_reg28_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg29 (
        .clk(comb_reg29_clk),
        .done(comb_reg29_done),
        .in(comb_reg29_in),
        .out(comb_reg29_out),
        .reset(comb_reg29_reset),
        .write_en(comb_reg29_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg30 (
        .clk(comb_reg30_clk),
        .done(comb_reg30_done),
        .in(comb_reg30_in),
        .out(comb_reg30_out),
        .reset(comb_reg30_reset),
        .write_en(comb_reg30_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) comb_reg31 (
        .clk(comb_reg31_clk),
        .done(comb_reg31_done),
        .in(comb_reg31_in),
        .out(comb_reg31_out),
        .reset(comb_reg31_reset),
        .write_en(comb_reg31_write_en)
    );
    std_reg # (
        .WIDTH(5)
    ) out (
        .clk(out_clk),
        .done(out_done),
        .in(out_in),
        .out(out_out),
        .reset(out_reset),
        .write_en(out_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm (
        .clk(fsm_clk),
        .done(fsm_done),
        .in(fsm_in),
        .out(fsm_out),
        .reset(fsm_reset),
        .write_en(fsm_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd (
        .clk(pd_clk),
        .done(pd_done),
        .in(pd_in),
        .out(pd_out),
        .reset(pd_reset),
        .write_en(pd_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm0 (
        .clk(fsm0_clk),
        .done(fsm0_done),
        .in(fsm0_in),
        .out(fsm0_out),
        .reset(fsm0_reset),
        .write_en(fsm0_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd0 (
        .clk(pd0_clk),
        .done(pd0_done),
        .in(pd0_in),
        .out(pd0_out),
        .reset(pd0_reset),
        .write_en(pd0_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm1 (
        .clk(fsm1_clk),
        .done(fsm1_done),
        .in(fsm1_in),
        .out(fsm1_out),
        .reset(fsm1_reset),
        .write_en(fsm1_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd1 (
        .clk(pd1_clk),
        .done(pd1_done),
        .in(pd1_in),
        .out(pd1_out),
        .reset(pd1_reset),
        .write_en(pd1_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm2 (
        .clk(fsm2_clk),
        .done(fsm2_done),
        .in(fsm2_in),
        .out(fsm2_out),
        .reset(fsm2_reset),
        .write_en(fsm2_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd2 (
        .clk(pd2_clk),
        .done(pd2_done),
        .in(pd2_in),
        .out(pd2_out),
        .reset(pd2_reset),
        .write_en(pd2_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm3 (
        .clk(fsm3_clk),
        .done(fsm3_done),
        .in(fsm3_in),
        .out(fsm3_out),
        .reset(fsm3_reset),
        .write_en(fsm3_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd3 (
        .clk(pd3_clk),
        .done(pd3_done),
        .in(pd3_in),
        .out(pd3_out),
        .reset(pd3_reset),
        .write_en(pd3_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm4 (
        .clk(fsm4_clk),
        .done(fsm4_done),
        .in(fsm4_in),
        .out(fsm4_out),
        .reset(fsm4_reset),
        .write_en(fsm4_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd4 (
        .clk(pd4_clk),
        .done(pd4_done),
        .in(pd4_in),
        .out(pd4_out),
        .reset(pd4_reset),
        .write_en(pd4_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm5 (
        .clk(fsm5_clk),
        .done(fsm5_done),
        .in(fsm5_in),
        .out(fsm5_out),
        .reset(fsm5_reset),
        .write_en(fsm5_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd5 (
        .clk(pd5_clk),
        .done(pd5_done),
        .in(pd5_in),
        .out(pd5_out),
        .reset(pd5_reset),
        .write_en(pd5_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm6 (
        .clk(fsm6_clk),
        .done(fsm6_done),
        .in(fsm6_in),
        .out(fsm6_out),
        .reset(fsm6_reset),
        .write_en(fsm6_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd6 (
        .clk(pd6_clk),
        .done(pd6_done),
        .in(pd6_in),
        .out(pd6_out),
        .reset(pd6_reset),
        .write_en(pd6_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm7 (
        .clk(fsm7_clk),
        .done(fsm7_done),
        .in(fsm7_in),
        .out(fsm7_out),
        .reset(fsm7_reset),
        .write_en(fsm7_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd7 (
        .clk(pd7_clk),
        .done(pd7_done),
        .in(pd7_in),
        .out(pd7_out),
        .reset(pd7_reset),
        .write_en(pd7_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm8 (
        .clk(fsm8_clk),
        .done(fsm8_done),
        .in(fsm8_in),
        .out(fsm8_out),
        .reset(fsm8_reset),
        .write_en(fsm8_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd8 (
        .clk(pd8_clk),
        .done(pd8_done),
        .in(pd8_in),
        .out(pd8_out),
        .reset(pd8_reset),
        .write_en(pd8_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm9 (
        .clk(fsm9_clk),
        .done(fsm9_done),
        .in(fsm9_in),
        .out(fsm9_out),
        .reset(fsm9_reset),
        .write_en(fsm9_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd9 (
        .clk(pd9_clk),
        .done(pd9_done),
        .in(pd9_in),
        .out(pd9_out),
        .reset(pd9_reset),
        .write_en(pd9_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm10 (
        .clk(fsm10_clk),
        .done(fsm10_done),
        .in(fsm10_in),
        .out(fsm10_out),
        .reset(fsm10_reset),
        .write_en(fsm10_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd10 (
        .clk(pd10_clk),
        .done(pd10_done),
        .in(pd10_in),
        .out(pd10_out),
        .reset(pd10_reset),
        .write_en(pd10_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm11 (
        .clk(fsm11_clk),
        .done(fsm11_done),
        .in(fsm11_in),
        .out(fsm11_out),
        .reset(fsm11_reset),
        .write_en(fsm11_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd11 (
        .clk(pd11_clk),
        .done(pd11_done),
        .in(pd11_in),
        .out(pd11_out),
        .reset(pd11_reset),
        .write_en(pd11_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm12 (
        .clk(fsm12_clk),
        .done(fsm12_done),
        .in(fsm12_in),
        .out(fsm12_out),
        .reset(fsm12_reset),
        .write_en(fsm12_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd12 (
        .clk(pd12_clk),
        .done(pd12_done),
        .in(pd12_in),
        .out(pd12_out),
        .reset(pd12_reset),
        .write_en(pd12_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm13 (
        .clk(fsm13_clk),
        .done(fsm13_done),
        .in(fsm13_in),
        .out(fsm13_out),
        .reset(fsm13_reset),
        .write_en(fsm13_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd13 (
        .clk(pd13_clk),
        .done(pd13_done),
        .in(pd13_in),
        .out(pd13_out),
        .reset(pd13_reset),
        .write_en(pd13_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm14 (
        .clk(fsm14_clk),
        .done(fsm14_done),
        .in(fsm14_in),
        .out(fsm14_out),
        .reset(fsm14_reset),
        .write_en(fsm14_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd14 (
        .clk(pd14_clk),
        .done(pd14_done),
        .in(pd14_in),
        .out(pd14_out),
        .reset(pd14_reset),
        .write_en(pd14_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm15 (
        .clk(fsm15_clk),
        .done(fsm15_done),
        .in(fsm15_in),
        .out(fsm15_out),
        .reset(fsm15_reset),
        .write_en(fsm15_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd15 (
        .clk(pd15_clk),
        .done(pd15_done),
        .in(pd15_in),
        .out(pd15_out),
        .reset(pd15_reset),
        .write_en(pd15_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm16 (
        .clk(fsm16_clk),
        .done(fsm16_done),
        .in(fsm16_in),
        .out(fsm16_out),
        .reset(fsm16_reset),
        .write_en(fsm16_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd16 (
        .clk(pd16_clk),
        .done(pd16_done),
        .in(pd16_in),
        .out(pd16_out),
        .reset(pd16_reset),
        .write_en(pd16_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm17 (
        .clk(fsm17_clk),
        .done(fsm17_done),
        .in(fsm17_in),
        .out(fsm17_out),
        .reset(fsm17_reset),
        .write_en(fsm17_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd17 (
        .clk(pd17_clk),
        .done(pd17_done),
        .in(pd17_in),
        .out(pd17_out),
        .reset(pd17_reset),
        .write_en(pd17_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm18 (
        .clk(fsm18_clk),
        .done(fsm18_done),
        .in(fsm18_in),
        .out(fsm18_out),
        .reset(fsm18_reset),
        .write_en(fsm18_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd18 (
        .clk(pd18_clk),
        .done(pd18_done),
        .in(pd18_in),
        .out(pd18_out),
        .reset(pd18_reset),
        .write_en(pd18_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm19 (
        .clk(fsm19_clk),
        .done(fsm19_done),
        .in(fsm19_in),
        .out(fsm19_out),
        .reset(fsm19_reset),
        .write_en(fsm19_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd19 (
        .clk(pd19_clk),
        .done(pd19_done),
        .in(pd19_in),
        .out(pd19_out),
        .reset(pd19_reset),
        .write_en(pd19_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm20 (
        .clk(fsm20_clk),
        .done(fsm20_done),
        .in(fsm20_in),
        .out(fsm20_out),
        .reset(fsm20_reset),
        .write_en(fsm20_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd20 (
        .clk(pd20_clk),
        .done(pd20_done),
        .in(pd20_in),
        .out(pd20_out),
        .reset(pd20_reset),
        .write_en(pd20_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm21 (
        .clk(fsm21_clk),
        .done(fsm21_done),
        .in(fsm21_in),
        .out(fsm21_out),
        .reset(fsm21_reset),
        .write_en(fsm21_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd21 (
        .clk(pd21_clk),
        .done(pd21_done),
        .in(pd21_in),
        .out(pd21_out),
        .reset(pd21_reset),
        .write_en(pd21_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm22 (
        .clk(fsm22_clk),
        .done(fsm22_done),
        .in(fsm22_in),
        .out(fsm22_out),
        .reset(fsm22_reset),
        .write_en(fsm22_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd22 (
        .clk(pd22_clk),
        .done(pd22_done),
        .in(pd22_in),
        .out(pd22_out),
        .reset(pd22_reset),
        .write_en(pd22_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm23 (
        .clk(fsm23_clk),
        .done(fsm23_done),
        .in(fsm23_in),
        .out(fsm23_out),
        .reset(fsm23_reset),
        .write_en(fsm23_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd23 (
        .clk(pd23_clk),
        .done(pd23_done),
        .in(pd23_in),
        .out(pd23_out),
        .reset(pd23_reset),
        .write_en(pd23_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm24 (
        .clk(fsm24_clk),
        .done(fsm24_done),
        .in(fsm24_in),
        .out(fsm24_out),
        .reset(fsm24_reset),
        .write_en(fsm24_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd24 (
        .clk(pd24_clk),
        .done(pd24_done),
        .in(pd24_in),
        .out(pd24_out),
        .reset(pd24_reset),
        .write_en(pd24_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm25 (
        .clk(fsm25_clk),
        .done(fsm25_done),
        .in(fsm25_in),
        .out(fsm25_out),
        .reset(fsm25_reset),
        .write_en(fsm25_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd25 (
        .clk(pd25_clk),
        .done(pd25_done),
        .in(pd25_in),
        .out(pd25_out),
        .reset(pd25_reset),
        .write_en(pd25_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm26 (
        .clk(fsm26_clk),
        .done(fsm26_done),
        .in(fsm26_in),
        .out(fsm26_out),
        .reset(fsm26_reset),
        .write_en(fsm26_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd26 (
        .clk(pd26_clk),
        .done(pd26_done),
        .in(pd26_in),
        .out(pd26_out),
        .reset(pd26_reset),
        .write_en(pd26_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm27 (
        .clk(fsm27_clk),
        .done(fsm27_done),
        .in(fsm27_in),
        .out(fsm27_out),
        .reset(fsm27_reset),
        .write_en(fsm27_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd27 (
        .clk(pd27_clk),
        .done(pd27_done),
        .in(pd27_in),
        .out(pd27_out),
        .reset(pd27_reset),
        .write_en(pd27_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm28 (
        .clk(fsm28_clk),
        .done(fsm28_done),
        .in(fsm28_in),
        .out(fsm28_out),
        .reset(fsm28_reset),
        .write_en(fsm28_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd28 (
        .clk(pd28_clk),
        .done(pd28_done),
        .in(pd28_in),
        .out(pd28_out),
        .reset(pd28_reset),
        .write_en(pd28_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm29 (
        .clk(fsm29_clk),
        .done(fsm29_done),
        .in(fsm29_in),
        .out(fsm29_out),
        .reset(fsm29_reset),
        .write_en(fsm29_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd29 (
        .clk(pd29_clk),
        .done(pd29_done),
        .in(pd29_in),
        .out(pd29_out),
        .reset(pd29_reset),
        .write_en(pd29_write_en)
    );
    std_reg # (
        .WIDTH(2)
    ) fsm30 (
        .clk(fsm30_clk),
        .done(fsm30_done),
        .in(fsm30_in),
        .out(fsm30_out),
        .reset(fsm30_reset),
        .write_en(fsm30_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd30 (
        .clk(pd30_clk),
        .done(pd30_done),
        .in(pd30_in),
        .out(pd30_out),
        .reset(pd30_reset),
        .write_en(pd30_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd31 (
        .clk(pd31_clk),
        .done(pd31_done),
        .in(pd31_in),
        .out(pd31_out),
        .reset(pd31_reset),
        .write_en(pd31_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd32 (
        .clk(pd32_clk),
        .done(pd32_done),
        .in(pd32_in),
        .out(pd32_out),
        .reset(pd32_reset),
        .write_en(pd32_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd33 (
        .clk(pd33_clk),
        .done(pd33_done),
        .in(pd33_in),
        .out(pd33_out),
        .reset(pd33_reset),
        .write_en(pd33_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd34 (
        .clk(pd34_clk),
        .done(pd34_done),
        .in(pd34_in),
        .out(pd34_out),
        .reset(pd34_reset),
        .write_en(pd34_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd35 (
        .clk(pd35_clk),
        .done(pd35_done),
        .in(pd35_in),
        .out(pd35_out),
        .reset(pd35_reset),
        .write_en(pd35_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd36 (
        .clk(pd36_clk),
        .done(pd36_done),
        .in(pd36_in),
        .out(pd36_out),
        .reset(pd36_reset),
        .write_en(pd36_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd37 (
        .clk(pd37_clk),
        .done(pd37_done),
        .in(pd37_in),
        .out(pd37_out),
        .reset(pd37_reset),
        .write_en(pd37_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd38 (
        .clk(pd38_clk),
        .done(pd38_done),
        .in(pd38_in),
        .out(pd38_out),
        .reset(pd38_reset),
        .write_en(pd38_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd39 (
        .clk(pd39_clk),
        .done(pd39_done),
        .in(pd39_in),
        .out(pd39_out),
        .reset(pd39_reset),
        .write_en(pd39_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd40 (
        .clk(pd40_clk),
        .done(pd40_done),
        .in(pd40_in),
        .out(pd40_out),
        .reset(pd40_reset),
        .write_en(pd40_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd41 (
        .clk(pd41_clk),
        .done(pd41_done),
        .in(pd41_in),
        .out(pd41_out),
        .reset(pd41_reset),
        .write_en(pd41_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd42 (
        .clk(pd42_clk),
        .done(pd42_done),
        .in(pd42_in),
        .out(pd42_out),
        .reset(pd42_reset),
        .write_en(pd42_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd43 (
        .clk(pd43_clk),
        .done(pd43_done),
        .in(pd43_in),
        .out(pd43_out),
        .reset(pd43_reset),
        .write_en(pd43_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd44 (
        .clk(pd44_clk),
        .done(pd44_done),
        .in(pd44_in),
        .out(pd44_out),
        .reset(pd44_reset),
        .write_en(pd44_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd45 (
        .clk(pd45_clk),
        .done(pd45_done),
        .in(pd45_in),
        .out(pd45_out),
        .reset(pd45_reset),
        .write_en(pd45_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd46 (
        .clk(pd46_clk),
        .done(pd46_done),
        .in(pd46_in),
        .out(pd46_out),
        .reset(pd46_reset),
        .write_en(pd46_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd47 (
        .clk(pd47_clk),
        .done(pd47_done),
        .in(pd47_in),
        .out(pd47_out),
        .reset(pd47_reset),
        .write_en(pd47_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd48 (
        .clk(pd48_clk),
        .done(pd48_done),
        .in(pd48_in),
        .out(pd48_out),
        .reset(pd48_reset),
        .write_en(pd48_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd49 (
        .clk(pd49_clk),
        .done(pd49_done),
        .in(pd49_in),
        .out(pd49_out),
        .reset(pd49_reset),
        .write_en(pd49_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd50 (
        .clk(pd50_clk),
        .done(pd50_done),
        .in(pd50_in),
        .out(pd50_out),
        .reset(pd50_reset),
        .write_en(pd50_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd51 (
        .clk(pd51_clk),
        .done(pd51_done),
        .in(pd51_in),
        .out(pd51_out),
        .reset(pd51_reset),
        .write_en(pd51_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd52 (
        .clk(pd52_clk),
        .done(pd52_done),
        .in(pd52_in),
        .out(pd52_out),
        .reset(pd52_reset),
        .write_en(pd52_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd53 (
        .clk(pd53_clk),
        .done(pd53_done),
        .in(pd53_in),
        .out(pd53_out),
        .reset(pd53_reset),
        .write_en(pd53_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd54 (
        .clk(pd54_clk),
        .done(pd54_done),
        .in(pd54_in),
        .out(pd54_out),
        .reset(pd54_reset),
        .write_en(pd54_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd55 (
        .clk(pd55_clk),
        .done(pd55_done),
        .in(pd55_in),
        .out(pd55_out),
        .reset(pd55_reset),
        .write_en(pd55_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd56 (
        .clk(pd56_clk),
        .done(pd56_done),
        .in(pd56_in),
        .out(pd56_out),
        .reset(pd56_reset),
        .write_en(pd56_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd57 (
        .clk(pd57_clk),
        .done(pd57_done),
        .in(pd57_in),
        .out(pd57_out),
        .reset(pd57_reset),
        .write_en(pd57_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd58 (
        .clk(pd58_clk),
        .done(pd58_done),
        .in(pd58_in),
        .out(pd58_out),
        .reset(pd58_reset),
        .write_en(pd58_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd59 (
        .clk(pd59_clk),
        .done(pd59_done),
        .in(pd59_in),
        .out(pd59_out),
        .reset(pd59_reset),
        .write_en(pd59_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd60 (
        .clk(pd60_clk),
        .done(pd60_done),
        .in(pd60_in),
        .out(pd60_out),
        .reset(pd60_reset),
        .write_en(pd60_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd61 (
        .clk(pd61_clk),
        .done(pd61_done),
        .in(pd61_in),
        .out(pd61_out),
        .reset(pd61_reset),
        .write_en(pd61_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd62 (
        .clk(pd62_clk),
        .done(pd62_done),
        .in(pd62_in),
        .out(pd62_out),
        .reset(pd62_reset),
        .write_en(pd62_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd63 (
        .clk(pd63_clk),
        .done(pd63_done),
        .in(pd63_in),
        .out(pd63_out),
        .reset(pd63_reset),
        .write_en(pd63_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd64 (
        .clk(pd64_clk),
        .done(pd64_done),
        .in(pd64_in),
        .out(pd64_out),
        .reset(pd64_reset),
        .write_en(pd64_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd65 (
        .clk(pd65_clk),
        .done(pd65_done),
        .in(pd65_in),
        .out(pd65_out),
        .reset(pd65_reset),
        .write_en(pd65_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd66 (
        .clk(pd66_clk),
        .done(pd66_done),
        .in(pd66_in),
        .out(pd66_out),
        .reset(pd66_reset),
        .write_en(pd66_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd67 (
        .clk(pd67_clk),
        .done(pd67_done),
        .in(pd67_in),
        .out(pd67_out),
        .reset(pd67_reset),
        .write_en(pd67_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd68 (
        .clk(pd68_clk),
        .done(pd68_done),
        .in(pd68_in),
        .out(pd68_out),
        .reset(pd68_reset),
        .write_en(pd68_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd69 (
        .clk(pd69_clk),
        .done(pd69_done),
        .in(pd69_in),
        .out(pd69_out),
        .reset(pd69_reset),
        .write_en(pd69_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd70 (
        .clk(pd70_clk),
        .done(pd70_done),
        .in(pd70_in),
        .out(pd70_out),
        .reset(pd70_reset),
        .write_en(pd70_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd71 (
        .clk(pd71_clk),
        .done(pd71_done),
        .in(pd71_in),
        .out(pd71_out),
        .reset(pd71_reset),
        .write_en(pd71_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd72 (
        .clk(pd72_clk),
        .done(pd72_done),
        .in(pd72_in),
        .out(pd72_out),
        .reset(pd72_reset),
        .write_en(pd72_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd73 (
        .clk(pd73_clk),
        .done(pd73_done),
        .in(pd73_in),
        .out(pd73_out),
        .reset(pd73_reset),
        .write_en(pd73_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd74 (
        .clk(pd74_clk),
        .done(pd74_done),
        .in(pd74_in),
        .out(pd74_out),
        .reset(pd74_reset),
        .write_en(pd74_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd75 (
        .clk(pd75_clk),
        .done(pd75_done),
        .in(pd75_in),
        .out(pd75_out),
        .reset(pd75_reset),
        .write_en(pd75_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd76 (
        .clk(pd76_clk),
        .done(pd76_done),
        .in(pd76_in),
        .out(pd76_out),
        .reset(pd76_reset),
        .write_en(pd76_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd77 (
        .clk(pd77_clk),
        .done(pd77_done),
        .in(pd77_in),
        .out(pd77_out),
        .reset(pd77_reset),
        .write_en(pd77_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd78 (
        .clk(pd78_clk),
        .done(pd78_done),
        .in(pd78_in),
        .out(pd78_out),
        .reset(pd78_reset),
        .write_en(pd78_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd79 (
        .clk(pd79_clk),
        .done(pd79_done),
        .in(pd79_in),
        .out(pd79_out),
        .reset(pd79_reset),
        .write_en(pd79_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd80 (
        .clk(pd80_clk),
        .done(pd80_done),
        .in(pd80_in),
        .out(pd80_out),
        .reset(pd80_reset),
        .write_en(pd80_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd81 (
        .clk(pd81_clk),
        .done(pd81_done),
        .in(pd81_in),
        .out(pd81_out),
        .reset(pd81_reset),
        .write_en(pd81_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd82 (
        .clk(pd82_clk),
        .done(pd82_done),
        .in(pd82_in),
        .out(pd82_out),
        .reset(pd82_reset),
        .write_en(pd82_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd83 (
        .clk(pd83_clk),
        .done(pd83_done),
        .in(pd83_in),
        .out(pd83_out),
        .reset(pd83_reset),
        .write_en(pd83_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd84 (
        .clk(pd84_clk),
        .done(pd84_done),
        .in(pd84_in),
        .out(pd84_out),
        .reset(pd84_reset),
        .write_en(pd84_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd85 (
        .clk(pd85_clk),
        .done(pd85_done),
        .in(pd85_in),
        .out(pd85_out),
        .reset(pd85_reset),
        .write_en(pd85_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd86 (
        .clk(pd86_clk),
        .done(pd86_done),
        .in(pd86_in),
        .out(pd86_out),
        .reset(pd86_reset),
        .write_en(pd86_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd87 (
        .clk(pd87_clk),
        .done(pd87_done),
        .in(pd87_in),
        .out(pd87_out),
        .reset(pd87_reset),
        .write_en(pd87_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd88 (
        .clk(pd88_clk),
        .done(pd88_done),
        .in(pd88_in),
        .out(pd88_out),
        .reset(pd88_reset),
        .write_en(pd88_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd89 (
        .clk(pd89_clk),
        .done(pd89_done),
        .in(pd89_in),
        .out(pd89_out),
        .reset(pd89_reset),
        .write_en(pd89_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd90 (
        .clk(pd90_clk),
        .done(pd90_done),
        .in(pd90_in),
        .out(pd90_out),
        .reset(pd90_reset),
        .write_en(pd90_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd91 (
        .clk(pd91_clk),
        .done(pd91_done),
        .in(pd91_in),
        .out(pd91_out),
        .reset(pd91_reset),
        .write_en(pd91_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd92 (
        .clk(pd92_clk),
        .done(pd92_done),
        .in(pd92_in),
        .out(pd92_out),
        .reset(pd92_reset),
        .write_en(pd92_write_en)
    );
    std_reg # (
        .WIDTH(3)
    ) fsm31 (
        .clk(fsm31_clk),
        .done(fsm31_done),
        .in(fsm31_in),
        .out(fsm31_out),
        .reset(fsm31_reset),
        .write_en(fsm31_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd93 (
        .clk(pd93_clk),
        .done(pd93_done),
        .in(pd93_in),
        .out(pd93_out),
        .reset(pd93_reset),
        .write_en(pd93_write_en)
    );
    std_reg # (
        .WIDTH(4)
    ) fsm32 (
        .clk(fsm32_clk),
        .done(fsm32_done),
        .in(fsm32_in),
        .out(fsm32_out),
        .reset(fsm32_reset),
        .write_en(fsm32_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) pd94 (
        .clk(pd94_clk),
        .done(pd94_done),
        .in(pd94_in),
        .out(pd94_out),
        .reset(pd94_reset),
        .write_en(pd94_write_en)
    );
    std_reg # (
        .WIDTH(1)
    ) fsm33 (
        .clk(fsm33_clk),
        .done(fsm33_done),
        .in(fsm33_in),
        .out(fsm33_out),
        .reset(fsm33_reset),
        .write_en(fsm33_write_en)
    );
    std_wire # (
        .WIDTH(1)
    ) write_zero_go (
        .in(write_zero_go_in),
        .out(write_zero_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write_zero_done (
        .in(write_zero_done_in),
        .out(write_zero_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write0_go (
        .in(write0_go_in),
        .out(write0_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write0_done (
        .in(write0_done_in),
        .out(write0_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write1_go (
        .in(write1_go_in),
        .out(write1_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write1_done (
        .in(write1_done_in),
        .out(write1_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write2_go (
        .in(write2_go_in),
        .out(write2_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write2_done (
        .in(write2_done_in),
        .out(write2_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write3_go (
        .in(write3_go_in),
        .out(write3_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write3_done (
        .in(write3_done_in),
        .out(write3_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write4_go (
        .in(write4_go_in),
        .out(write4_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write4_done (
        .in(write4_done_in),
        .out(write4_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write5_go (
        .in(write5_go_in),
        .out(write5_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write5_done (
        .in(write5_done_in),
        .out(write5_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write6_go (
        .in(write6_go_in),
        .out(write6_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write6_done (
        .in(write6_done_in),
        .out(write6_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write7_go (
        .in(write7_go_in),
        .out(write7_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write7_done (
        .in(write7_done_in),
        .out(write7_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write8_go (
        .in(write8_go_in),
        .out(write8_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write8_done (
        .in(write8_done_in),
        .out(write8_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write9_go (
        .in(write9_go_in),
        .out(write9_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write9_done (
        .in(write9_done_in),
        .out(write9_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write10_go (
        .in(write10_go_in),
        .out(write10_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write10_done (
        .in(write10_done_in),
        .out(write10_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write11_go (
        .in(write11_go_in),
        .out(write11_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write11_done (
        .in(write11_done_in),
        .out(write11_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write12_go (
        .in(write12_go_in),
        .out(write12_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write12_done (
        .in(write12_done_in),
        .out(write12_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write13_go (
        .in(write13_go_in),
        .out(write13_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write13_done (
        .in(write13_done_in),
        .out(write13_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write14_go (
        .in(write14_go_in),
        .out(write14_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write14_done (
        .in(write14_done_in),
        .out(write14_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write15_go (
        .in(write15_go_in),
        .out(write15_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write15_done (
        .in(write15_done_in),
        .out(write15_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write16_go (
        .in(write16_go_in),
        .out(write16_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write16_done (
        .in(write16_done_in),
        .out(write16_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write17_go (
        .in(write17_go_in),
        .out(write17_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write17_done (
        .in(write17_done_in),
        .out(write17_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write18_go (
        .in(write18_go_in),
        .out(write18_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write18_done (
        .in(write18_done_in),
        .out(write18_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write19_go (
        .in(write19_go_in),
        .out(write19_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write19_done (
        .in(write19_done_in),
        .out(write19_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write20_go (
        .in(write20_go_in),
        .out(write20_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write20_done (
        .in(write20_done_in),
        .out(write20_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write21_go (
        .in(write21_go_in),
        .out(write21_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write21_done (
        .in(write21_done_in),
        .out(write21_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write22_go (
        .in(write22_go_in),
        .out(write22_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write22_done (
        .in(write22_done_in),
        .out(write22_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write23_go (
        .in(write23_go_in),
        .out(write23_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write23_done (
        .in(write23_done_in),
        .out(write23_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write24_go (
        .in(write24_go_in),
        .out(write24_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write24_done (
        .in(write24_done_in),
        .out(write24_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write25_go (
        .in(write25_go_in),
        .out(write25_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write25_done (
        .in(write25_done_in),
        .out(write25_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write26_go (
        .in(write26_go_in),
        .out(write26_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write26_done (
        .in(write26_done_in),
        .out(write26_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write27_go (
        .in(write27_go_in),
        .out(write27_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write27_done (
        .in(write27_done_in),
        .out(write27_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write28_go (
        .in(write28_go_in),
        .out(write28_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write28_done (
        .in(write28_done_in),
        .out(write28_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write29_go (
        .in(write29_go_in),
        .out(write29_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write29_done (
        .in(write29_done_in),
        .out(write29_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write30_go (
        .in(write30_go_in),
        .out(write30_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write30_done (
        .in(write30_done_in),
        .out(write30_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write31_go (
        .in(write31_go_in),
        .out(write31_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) write31_done (
        .in(write31_done_in),
        .out(write31_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) find_write_index_go (
        .in(find_write_index_go_in),
        .out(find_write_index_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) find_write_index_done (
        .in(find_write_index_done_in),
        .out(find_write_index_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) default_to_zero_length_index_go (
        .in(default_to_zero_length_index_go_in),
        .out(default_to_zero_length_index_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) default_to_zero_length_index_done (
        .in(default_to_zero_length_index_done_in),
        .out(default_to_zero_length_index_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) save_index_go (
        .in(save_index_go_in),
        .out(save_index_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) save_index_done (
        .in(save_index_done_in),
        .out(save_index_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) is_length_zero0_go (
        .in(is_length_zero0_go_in),
        .out(is_length_zero0_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) is_length_zero0_done (
        .in(is_length_zero0_done_in),
        .out(is_length_zero0_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke_go (
        .in(invoke_go_in),
        .out(invoke_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke_done (
        .in(invoke_done_in),
        .out(invoke_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke0_go (
        .in(invoke0_go_in),
        .out(invoke0_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke0_done (
        .in(invoke0_done_in),
        .out(invoke0_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke1_go (
        .in(invoke1_go_in),
        .out(invoke1_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke1_done (
        .in(invoke1_done_in),
        .out(invoke1_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke2_go (
        .in(invoke2_go_in),
        .out(invoke2_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke2_done (
        .in(invoke2_done_in),
        .out(invoke2_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke3_go (
        .in(invoke3_go_in),
        .out(invoke3_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke3_done (
        .in(invoke3_done_in),
        .out(invoke3_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke4_go (
        .in(invoke4_go_in),
        .out(invoke4_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke4_done (
        .in(invoke4_done_in),
        .out(invoke4_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke5_go (
        .in(invoke5_go_in),
        .out(invoke5_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke5_done (
        .in(invoke5_done_in),
        .out(invoke5_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke6_go (
        .in(invoke6_go_in),
        .out(invoke6_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke6_done (
        .in(invoke6_done_in),
        .out(invoke6_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke7_go (
        .in(invoke7_go_in),
        .out(invoke7_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke7_done (
        .in(invoke7_done_in),
        .out(invoke7_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke8_go (
        .in(invoke8_go_in),
        .out(invoke8_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke8_done (
        .in(invoke8_done_in),
        .out(invoke8_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke9_go (
        .in(invoke9_go_in),
        .out(invoke9_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke9_done (
        .in(invoke9_done_in),
        .out(invoke9_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke10_go (
        .in(invoke10_go_in),
        .out(invoke10_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke10_done (
        .in(invoke10_done_in),
        .out(invoke10_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke11_go (
        .in(invoke11_go_in),
        .out(invoke11_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke11_done (
        .in(invoke11_done_in),
        .out(invoke11_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke12_go (
        .in(invoke12_go_in),
        .out(invoke12_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke12_done (
        .in(invoke12_done_in),
        .out(invoke12_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke13_go (
        .in(invoke13_go_in),
        .out(invoke13_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke13_done (
        .in(invoke13_done_in),
        .out(invoke13_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke14_go (
        .in(invoke14_go_in),
        .out(invoke14_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke14_done (
        .in(invoke14_done_in),
        .out(invoke14_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke15_go (
        .in(invoke15_go_in),
        .out(invoke15_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke15_done (
        .in(invoke15_done_in),
        .out(invoke15_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke16_go (
        .in(invoke16_go_in),
        .out(invoke16_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke16_done (
        .in(invoke16_done_in),
        .out(invoke16_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke17_go (
        .in(invoke17_go_in),
        .out(invoke17_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke17_done (
        .in(invoke17_done_in),
        .out(invoke17_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke18_go (
        .in(invoke18_go_in),
        .out(invoke18_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke18_done (
        .in(invoke18_done_in),
        .out(invoke18_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke19_go (
        .in(invoke19_go_in),
        .out(invoke19_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke19_done (
        .in(invoke19_done_in),
        .out(invoke19_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke20_go (
        .in(invoke20_go_in),
        .out(invoke20_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke20_done (
        .in(invoke20_done_in),
        .out(invoke20_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke21_go (
        .in(invoke21_go_in),
        .out(invoke21_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke21_done (
        .in(invoke21_done_in),
        .out(invoke21_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke22_go (
        .in(invoke22_go_in),
        .out(invoke22_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke22_done (
        .in(invoke22_done_in),
        .out(invoke22_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke23_go (
        .in(invoke23_go_in),
        .out(invoke23_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke23_done (
        .in(invoke23_done_in),
        .out(invoke23_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke24_go (
        .in(invoke24_go_in),
        .out(invoke24_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke24_done (
        .in(invoke24_done_in),
        .out(invoke24_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke25_go (
        .in(invoke25_go_in),
        .out(invoke25_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke25_done (
        .in(invoke25_done_in),
        .out(invoke25_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke26_go (
        .in(invoke26_go_in),
        .out(invoke26_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke26_done (
        .in(invoke26_done_in),
        .out(invoke26_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke27_go (
        .in(invoke27_go_in),
        .out(invoke27_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke27_done (
        .in(invoke27_done_in),
        .out(invoke27_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke28_go (
        .in(invoke28_go_in),
        .out(invoke28_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke28_done (
        .in(invoke28_done_in),
        .out(invoke28_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke29_go (
        .in(invoke29_go_in),
        .out(invoke29_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke29_done (
        .in(invoke29_done_in),
        .out(invoke29_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke30_go (
        .in(invoke30_go_in),
        .out(invoke30_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke30_done (
        .in(invoke30_done_in),
        .out(invoke30_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke31_go (
        .in(invoke31_go_in),
        .out(invoke31_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke31_done (
        .in(invoke31_done_in),
        .out(invoke31_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke32_go (
        .in(invoke32_go_in),
        .out(invoke32_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke32_done (
        .in(invoke32_done_in),
        .out(invoke32_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke33_go (
        .in(invoke33_go_in),
        .out(invoke33_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke33_done (
        .in(invoke33_done_in),
        .out(invoke33_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke34_go (
        .in(invoke34_go_in),
        .out(invoke34_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke34_done (
        .in(invoke34_done_in),
        .out(invoke34_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke35_go (
        .in(invoke35_go_in),
        .out(invoke35_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke35_done (
        .in(invoke35_done_in),
        .out(invoke35_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke36_go (
        .in(invoke36_go_in),
        .out(invoke36_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke36_done (
        .in(invoke36_done_in),
        .out(invoke36_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke37_go (
        .in(invoke37_go_in),
        .out(invoke37_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke37_done (
        .in(invoke37_done_in),
        .out(invoke37_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke38_go (
        .in(invoke38_go_in),
        .out(invoke38_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke38_done (
        .in(invoke38_done_in),
        .out(invoke38_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke39_go (
        .in(invoke39_go_in),
        .out(invoke39_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke39_done (
        .in(invoke39_done_in),
        .out(invoke39_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke40_go (
        .in(invoke40_go_in),
        .out(invoke40_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke40_done (
        .in(invoke40_done_in),
        .out(invoke40_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke41_go (
        .in(invoke41_go_in),
        .out(invoke41_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke41_done (
        .in(invoke41_done_in),
        .out(invoke41_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke42_go (
        .in(invoke42_go_in),
        .out(invoke42_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke42_done (
        .in(invoke42_done_in),
        .out(invoke42_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke43_go (
        .in(invoke43_go_in),
        .out(invoke43_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke43_done (
        .in(invoke43_done_in),
        .out(invoke43_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke44_go (
        .in(invoke44_go_in),
        .out(invoke44_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke44_done (
        .in(invoke44_done_in),
        .out(invoke44_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke45_go (
        .in(invoke45_go_in),
        .out(invoke45_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke45_done (
        .in(invoke45_done_in),
        .out(invoke45_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke46_go (
        .in(invoke46_go_in),
        .out(invoke46_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke46_done (
        .in(invoke46_done_in),
        .out(invoke46_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke47_go (
        .in(invoke47_go_in),
        .out(invoke47_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke47_done (
        .in(invoke47_done_in),
        .out(invoke47_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke48_go (
        .in(invoke48_go_in),
        .out(invoke48_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke48_done (
        .in(invoke48_done_in),
        .out(invoke48_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke49_go (
        .in(invoke49_go_in),
        .out(invoke49_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke49_done (
        .in(invoke49_done_in),
        .out(invoke49_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke50_go (
        .in(invoke50_go_in),
        .out(invoke50_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke50_done (
        .in(invoke50_done_in),
        .out(invoke50_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke51_go (
        .in(invoke51_go_in),
        .out(invoke51_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke51_done (
        .in(invoke51_done_in),
        .out(invoke51_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke52_go (
        .in(invoke52_go_in),
        .out(invoke52_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke52_done (
        .in(invoke52_done_in),
        .out(invoke52_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke53_go (
        .in(invoke53_go_in),
        .out(invoke53_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke53_done (
        .in(invoke53_done_in),
        .out(invoke53_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke54_go (
        .in(invoke54_go_in),
        .out(invoke54_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke54_done (
        .in(invoke54_done_in),
        .out(invoke54_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke55_go (
        .in(invoke55_go_in),
        .out(invoke55_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke55_done (
        .in(invoke55_done_in),
        .out(invoke55_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke56_go (
        .in(invoke56_go_in),
        .out(invoke56_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke56_done (
        .in(invoke56_done_in),
        .out(invoke56_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke57_go (
        .in(invoke57_go_in),
        .out(invoke57_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke57_done (
        .in(invoke57_done_in),
        .out(invoke57_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke58_go (
        .in(invoke58_go_in),
        .out(invoke58_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke58_done (
        .in(invoke58_done_in),
        .out(invoke58_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke59_go (
        .in(invoke59_go_in),
        .out(invoke59_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke59_done (
        .in(invoke59_done_in),
        .out(invoke59_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke60_go (
        .in(invoke60_go_in),
        .out(invoke60_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke60_done (
        .in(invoke60_done_in),
        .out(invoke60_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke61_go (
        .in(invoke61_go_in),
        .out(invoke61_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) invoke61_done (
        .in(invoke61_done_in),
        .out(invoke61_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par_go (
        .in(par_go_in),
        .out(par_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par_done (
        .in(par_done_in),
        .out(par_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc_go (
        .in(tdcc_go_in),
        .out(tdcc_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc_done (
        .in(tdcc_done_in),
        .out(tdcc_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc0_go (
        .in(tdcc0_go_in),
        .out(tdcc0_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc0_done (
        .in(tdcc0_done_in),
        .out(tdcc0_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc1_go (
        .in(tdcc1_go_in),
        .out(tdcc1_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc1_done (
        .in(tdcc1_done_in),
        .out(tdcc1_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc2_go (
        .in(tdcc2_go_in),
        .out(tdcc2_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc2_done (
        .in(tdcc2_done_in),
        .out(tdcc2_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc3_go (
        .in(tdcc3_go_in),
        .out(tdcc3_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc3_done (
        .in(tdcc3_done_in),
        .out(tdcc3_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc4_go (
        .in(tdcc4_go_in),
        .out(tdcc4_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc4_done (
        .in(tdcc4_done_in),
        .out(tdcc4_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc5_go (
        .in(tdcc5_go_in),
        .out(tdcc5_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc5_done (
        .in(tdcc5_done_in),
        .out(tdcc5_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc6_go (
        .in(tdcc6_go_in),
        .out(tdcc6_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc6_done (
        .in(tdcc6_done_in),
        .out(tdcc6_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc7_go (
        .in(tdcc7_go_in),
        .out(tdcc7_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc7_done (
        .in(tdcc7_done_in),
        .out(tdcc7_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc8_go (
        .in(tdcc8_go_in),
        .out(tdcc8_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc8_done (
        .in(tdcc8_done_in),
        .out(tdcc8_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc9_go (
        .in(tdcc9_go_in),
        .out(tdcc9_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc9_done (
        .in(tdcc9_done_in),
        .out(tdcc9_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc10_go (
        .in(tdcc10_go_in),
        .out(tdcc10_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc10_done (
        .in(tdcc10_done_in),
        .out(tdcc10_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc11_go (
        .in(tdcc11_go_in),
        .out(tdcc11_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc11_done (
        .in(tdcc11_done_in),
        .out(tdcc11_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc12_go (
        .in(tdcc12_go_in),
        .out(tdcc12_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc12_done (
        .in(tdcc12_done_in),
        .out(tdcc12_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc13_go (
        .in(tdcc13_go_in),
        .out(tdcc13_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc13_done (
        .in(tdcc13_done_in),
        .out(tdcc13_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc14_go (
        .in(tdcc14_go_in),
        .out(tdcc14_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc14_done (
        .in(tdcc14_done_in),
        .out(tdcc14_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc15_go (
        .in(tdcc15_go_in),
        .out(tdcc15_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc15_done (
        .in(tdcc15_done_in),
        .out(tdcc15_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc16_go (
        .in(tdcc16_go_in),
        .out(tdcc16_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc16_done (
        .in(tdcc16_done_in),
        .out(tdcc16_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc17_go (
        .in(tdcc17_go_in),
        .out(tdcc17_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc17_done (
        .in(tdcc17_done_in),
        .out(tdcc17_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc18_go (
        .in(tdcc18_go_in),
        .out(tdcc18_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc18_done (
        .in(tdcc18_done_in),
        .out(tdcc18_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc19_go (
        .in(tdcc19_go_in),
        .out(tdcc19_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc19_done (
        .in(tdcc19_done_in),
        .out(tdcc19_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc20_go (
        .in(tdcc20_go_in),
        .out(tdcc20_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc20_done (
        .in(tdcc20_done_in),
        .out(tdcc20_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc21_go (
        .in(tdcc21_go_in),
        .out(tdcc21_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc21_done (
        .in(tdcc21_done_in),
        .out(tdcc21_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc22_go (
        .in(tdcc22_go_in),
        .out(tdcc22_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc22_done (
        .in(tdcc22_done_in),
        .out(tdcc22_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc23_go (
        .in(tdcc23_go_in),
        .out(tdcc23_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc23_done (
        .in(tdcc23_done_in),
        .out(tdcc23_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc24_go (
        .in(tdcc24_go_in),
        .out(tdcc24_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc24_done (
        .in(tdcc24_done_in),
        .out(tdcc24_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc25_go (
        .in(tdcc25_go_in),
        .out(tdcc25_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc25_done (
        .in(tdcc25_done_in),
        .out(tdcc25_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc26_go (
        .in(tdcc26_go_in),
        .out(tdcc26_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc26_done (
        .in(tdcc26_done_in),
        .out(tdcc26_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc27_go (
        .in(tdcc27_go_in),
        .out(tdcc27_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc27_done (
        .in(tdcc27_done_in),
        .out(tdcc27_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc28_go (
        .in(tdcc28_go_in),
        .out(tdcc28_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc28_done (
        .in(tdcc28_done_in),
        .out(tdcc28_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc29_go (
        .in(tdcc29_go_in),
        .out(tdcc29_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc29_done (
        .in(tdcc29_done_in),
        .out(tdcc29_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc30_go (
        .in(tdcc30_go_in),
        .out(tdcc30_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc30_done (
        .in(tdcc30_done_in),
        .out(tdcc30_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par0_go (
        .in(par0_go_in),
        .out(par0_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par0_done (
        .in(par0_done_in),
        .out(par0_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par1_go (
        .in(par1_go_in),
        .out(par1_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par1_done (
        .in(par1_done_in),
        .out(par1_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par2_go (
        .in(par2_go_in),
        .out(par2_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par2_done (
        .in(par2_done_in),
        .out(par2_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par3_go (
        .in(par3_go_in),
        .out(par3_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par3_done (
        .in(par3_done_in),
        .out(par3_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par4_go (
        .in(par4_go_in),
        .out(par4_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par4_done (
        .in(par4_done_in),
        .out(par4_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par5_go (
        .in(par5_go_in),
        .out(par5_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) par5_done (
        .in(par5_done_in),
        .out(par5_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc31_go (
        .in(tdcc31_go_in),
        .out(tdcc31_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc31_done (
        .in(tdcc31_done_in),
        .out(tdcc31_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc32_go (
        .in(tdcc32_go_in),
        .out(tdcc32_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc32_done (
        .in(tdcc32_done_in),
        .out(tdcc32_done_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc33_go (
        .in(tdcc33_go_in),
        .out(tdcc33_go_out)
    );
    std_wire # (
        .WIDTH(1)
    ) tdcc33_done (
        .in(tdcc33_done_in),
        .out(tdcc33_done_out)
    );
    assign done = tdcc33_done_out;
    assign index = out_out;
    assign ce00_addrA =
     invoke31_go_out ? 5'd0 : 5'd0;
    assign ce00_addrB =
     invoke31_go_out ? 5'd1 : 5'd0;
    assign ce00_clk = clk;
    assign ce00_go = invoke31_go_out;
    assign ce00_lenA =
     invoke31_go_out ? l0_out : 5'd0;
    assign ce00_lenB =
     invoke31_go_out ? l1_out : 5'd0;
    assign ce00_mlA =
     invoke31_go_out ? me0_out : 1'd0;
    assign ce00_mlB =
     invoke31_go_out ? me1_out : 1'd0;
    assign ce00_reset = reset;
    assign ce01_addrA =
     invoke32_go_out ? 5'd2 : 5'd0;
    assign ce01_addrB =
     invoke32_go_out ? 5'd3 : 5'd0;
    assign ce01_clk = clk;
    assign ce01_go = invoke32_go_out;
    assign ce01_lenA =
     invoke32_go_out ? l2_out : 5'd0;
    assign ce01_lenB =
     invoke32_go_out ? l3_out : 5'd0;
    assign ce01_mlA =
     invoke32_go_out ? me2_out : 1'd0;
    assign ce01_mlB =
     invoke32_go_out ? me3_out : 1'd0;
    assign ce01_reset = reset;
    assign ce010_addrA =
     invoke41_go_out ? 5'd20 : 5'd0;
    assign ce010_addrB =
     invoke41_go_out ? 5'd21 : 5'd0;
    assign ce010_clk = clk;
    assign ce010_go = invoke41_go_out;
    assign ce010_lenA =
     invoke41_go_out ? l20_out : 5'd0;
    assign ce010_lenB =
     invoke41_go_out ? l21_out : 5'd0;
    assign ce010_mlA =
     invoke41_go_out ? me20_out : 1'd0;
    assign ce010_mlB =
     invoke41_go_out ? me21_out : 1'd0;
    assign ce010_reset = reset;
    assign ce011_addrA =
     invoke42_go_out ? 5'd22 : 5'd0;
    assign ce011_addrB =
     invoke42_go_out ? 5'd23 : 5'd0;
    assign ce011_clk = clk;
    assign ce011_go = invoke42_go_out;
    assign ce011_lenA =
     invoke42_go_out ? l22_out : 5'd0;
    assign ce011_lenB =
     invoke42_go_out ? l23_out : 5'd0;
    assign ce011_mlA =
     invoke42_go_out ? me22_out : 1'd0;
    assign ce011_mlB =
     invoke42_go_out ? me23_out : 1'd0;
    assign ce011_reset = reset;
    assign ce012_addrA =
     invoke43_go_out ? 5'd24 : 5'd0;
    assign ce012_addrB =
     invoke43_go_out ? 5'd25 : 5'd0;
    assign ce012_clk = clk;
    assign ce012_go = invoke43_go_out;
    assign ce012_lenA =
     invoke43_go_out ? l24_out : 5'd0;
    assign ce012_lenB =
     invoke43_go_out ? l25_out : 5'd0;
    assign ce012_mlA =
     invoke43_go_out ? me24_out : 1'd0;
    assign ce012_mlB =
     invoke43_go_out ? me25_out : 1'd0;
    assign ce012_reset = reset;
    assign ce013_addrA =
     invoke44_go_out ? 5'd26 : 5'd0;
    assign ce013_addrB =
     invoke44_go_out ? 5'd27 : 5'd0;
    assign ce013_clk = clk;
    assign ce013_go = invoke44_go_out;
    assign ce013_lenA =
     invoke44_go_out ? l26_out : 5'd0;
    assign ce013_lenB =
     invoke44_go_out ? l27_out : 5'd0;
    assign ce013_mlA =
     invoke44_go_out ? me26_out : 1'd0;
    assign ce013_mlB =
     invoke44_go_out ? me27_out : 1'd0;
    assign ce013_reset = reset;
    assign ce014_addrA =
     invoke45_go_out ? 5'd28 : 5'd0;
    assign ce014_addrB =
     invoke45_go_out ? 5'd29 : 5'd0;
    assign ce014_clk = clk;
    assign ce014_go = invoke45_go_out;
    assign ce014_lenA =
     invoke45_go_out ? l28_out : 5'd0;
    assign ce014_lenB =
     invoke45_go_out ? l29_out : 5'd0;
    assign ce014_mlA =
     invoke45_go_out ? me28_out : 1'd0;
    assign ce014_mlB =
     invoke45_go_out ? me29_out : 1'd0;
    assign ce014_reset = reset;
    assign ce015_addrA =
     invoke46_go_out ? 5'd30 : 5'd0;
    assign ce015_addrB =
     invoke46_go_out ? 5'd31 : 5'd0;
    assign ce015_clk = clk;
    assign ce015_go = invoke46_go_out;
    assign ce015_lenA =
     invoke46_go_out ? l30_out : 5'd0;
    assign ce015_lenB =
     invoke46_go_out ? l31_out : 5'd0;
    assign ce015_mlA =
     invoke46_go_out ? me30_out : 1'd0;
    assign ce015_mlB =
     invoke46_go_out ? me31_out : 1'd0;
    assign ce015_reset = reset;
    assign ce02_addrA =
     invoke33_go_out ? 5'd4 : 5'd0;
    assign ce02_addrB =
     invoke33_go_out ? 5'd5 : 5'd0;
    assign ce02_clk = clk;
    assign ce02_go = invoke33_go_out;
    assign ce02_lenA =
     invoke33_go_out ? l4_out : 5'd0;
    assign ce02_lenB =
     invoke33_go_out ? l5_out : 5'd0;
    assign ce02_mlA =
     invoke33_go_out ? me4_out : 1'd0;
    assign ce02_mlB =
     invoke33_go_out ? me5_out : 1'd0;
    assign ce02_reset = reset;
    assign ce03_addrA =
     invoke34_go_out ? 5'd6 : 5'd0;
    assign ce03_addrB =
     invoke34_go_out ? 5'd7 : 5'd0;
    assign ce03_clk = clk;
    assign ce03_go = invoke34_go_out;
    assign ce03_lenA =
     invoke34_go_out ? l6_out : 5'd0;
    assign ce03_lenB =
     invoke34_go_out ? l7_out : 5'd0;
    assign ce03_mlA =
     invoke34_go_out ? me6_out : 1'd0;
    assign ce03_mlB =
     invoke34_go_out ? me7_out : 1'd0;
    assign ce03_reset = reset;
    assign ce04_addrA =
     invoke35_go_out ? 5'd8 : 5'd0;
    assign ce04_addrB =
     invoke35_go_out ? 5'd9 : 5'd0;
    assign ce04_clk = clk;
    assign ce04_go = invoke35_go_out;
    assign ce04_lenA =
     invoke35_go_out ? l8_out : 5'd0;
    assign ce04_lenB =
     invoke35_go_out ? l9_out : 5'd0;
    assign ce04_mlA =
     invoke35_go_out ? me8_out : 1'd0;
    assign ce04_mlB =
     invoke35_go_out ? me9_out : 1'd0;
    assign ce04_reset = reset;
    assign ce05_addrA =
     invoke36_go_out ? 5'd10 : 5'd0;
    assign ce05_addrB =
     invoke36_go_out ? 5'd11 : 5'd0;
    assign ce05_clk = clk;
    assign ce05_go = invoke36_go_out;
    assign ce05_lenA =
     invoke36_go_out ? l10_out : 5'd0;
    assign ce05_lenB =
     invoke36_go_out ? l11_out : 5'd0;
    assign ce05_mlA =
     invoke36_go_out ? me10_out : 1'd0;
    assign ce05_mlB =
     invoke36_go_out ? me11_out : 1'd0;
    assign ce05_reset = reset;
    assign ce06_addrA =
     invoke37_go_out ? 5'd12 : 5'd0;
    assign ce06_addrB =
     invoke37_go_out ? 5'd13 : 5'd0;
    assign ce06_clk = clk;
    assign ce06_go = invoke37_go_out;
    assign ce06_lenA =
     invoke37_go_out ? l12_out : 5'd0;
    assign ce06_lenB =
     invoke37_go_out ? l13_out : 5'd0;
    assign ce06_mlA =
     invoke37_go_out ? me12_out : 1'd0;
    assign ce06_mlB =
     invoke37_go_out ? me13_out : 1'd0;
    assign ce06_reset = reset;
    assign ce07_addrA =
     invoke38_go_out ? 5'd14 : 5'd0;
    assign ce07_addrB =
     invoke38_go_out ? 5'd15 : 5'd0;
    assign ce07_clk = clk;
    assign ce07_go = invoke38_go_out;
    assign ce07_lenA =
     invoke38_go_out ? l14_out : 5'd0;
    assign ce07_lenB =
     invoke38_go_out ? l15_out : 5'd0;
    assign ce07_mlA =
     invoke38_go_out ? me14_out : 1'd0;
    assign ce07_mlB =
     invoke38_go_out ? me15_out : 1'd0;
    assign ce07_reset = reset;
    assign ce08_addrA =
     invoke39_go_out ? 5'd16 : 5'd0;
    assign ce08_addrB =
     invoke39_go_out ? 5'd17 : 5'd0;
    assign ce08_clk = clk;
    assign ce08_go = invoke39_go_out;
    assign ce08_lenA =
     invoke39_go_out ? l16_out : 5'd0;
    assign ce08_lenB =
     invoke39_go_out ? l17_out : 5'd0;
    assign ce08_mlA =
     invoke39_go_out ? me16_out : 1'd0;
    assign ce08_mlB =
     invoke39_go_out ? me17_out : 1'd0;
    assign ce08_reset = reset;
    assign ce09_addrA =
     invoke40_go_out ? 5'd18 : 5'd0;
    assign ce09_addrB =
     invoke40_go_out ? 5'd19 : 5'd0;
    assign ce09_clk = clk;
    assign ce09_go = invoke40_go_out;
    assign ce09_lenA =
     invoke40_go_out ? l18_out : 5'd0;
    assign ce09_lenB =
     invoke40_go_out ? l19_out : 5'd0;
    assign ce09_mlA =
     invoke40_go_out ? me18_out : 1'd0;
    assign ce09_mlB =
     invoke40_go_out ? me19_out : 1'd0;
    assign ce09_reset = reset;
    assign ce10_addrA =
     invoke47_go_out ? ce00_addrX : 5'd0;
    assign ce10_addrB =
     invoke47_go_out ? ce01_addrX : 5'd0;
    assign ce10_clk = clk;
    assign ce10_go = invoke47_go_out;
    assign ce10_lenA =
     invoke47_go_out ? ce00_lenX : 5'd0;
    assign ce10_lenB =
     invoke47_go_out ? ce01_lenX : 5'd0;
    assign ce10_mlA =
     invoke47_go_out ? ce00_mlX : 1'd0;
    assign ce10_mlB =
     invoke47_go_out ? ce01_mlX : 1'd0;
    assign ce10_reset = reset;
    assign ce11_addrA =
     invoke48_go_out ? ce02_addrX : 5'd0;
    assign ce11_addrB =
     invoke48_go_out ? ce03_addrX : 5'd0;
    assign ce11_clk = clk;
    assign ce11_go = invoke48_go_out;
    assign ce11_lenA =
     invoke48_go_out ? ce02_lenX : 5'd0;
    assign ce11_lenB =
     invoke48_go_out ? ce03_lenX : 5'd0;
    assign ce11_mlA =
     invoke48_go_out ? ce02_mlX : 1'd0;
    assign ce11_mlB =
     invoke48_go_out ? ce03_mlX : 1'd0;
    assign ce11_reset = reset;
    assign ce12_addrA =
     invoke49_go_out ? ce04_addrX : 5'd0;
    assign ce12_addrB =
     invoke49_go_out ? ce05_addrX : 5'd0;
    assign ce12_clk = clk;
    assign ce12_go = invoke49_go_out;
    assign ce12_lenA =
     invoke49_go_out ? ce04_lenX : 5'd0;
    assign ce12_lenB =
     invoke49_go_out ? ce05_lenX : 5'd0;
    assign ce12_mlA =
     invoke49_go_out ? ce04_mlX : 1'd0;
    assign ce12_mlB =
     invoke49_go_out ? ce05_mlX : 1'd0;
    assign ce12_reset = reset;
    assign ce13_addrA =
     invoke50_go_out ? ce06_addrX : 5'd0;
    assign ce13_addrB =
     invoke50_go_out ? ce07_addrX : 5'd0;
    assign ce13_clk = clk;
    assign ce13_go = invoke50_go_out;
    assign ce13_lenA =
     invoke50_go_out ? ce06_lenX : 5'd0;
    assign ce13_lenB =
     invoke50_go_out ? ce07_lenX : 5'd0;
    assign ce13_mlA =
     invoke50_go_out ? ce06_mlX : 1'd0;
    assign ce13_mlB =
     invoke50_go_out ? ce07_mlX : 1'd0;
    assign ce13_reset = reset;
    assign ce14_addrA =
     invoke51_go_out ? ce08_addrX : 5'd0;
    assign ce14_addrB =
     invoke51_go_out ? ce09_addrX : 5'd0;
    assign ce14_clk = clk;
    assign ce14_go = invoke51_go_out;
    assign ce14_lenA =
     invoke51_go_out ? ce08_lenX : 5'd0;
    assign ce14_lenB =
     invoke51_go_out ? ce09_lenX : 5'd0;
    assign ce14_mlA =
     invoke51_go_out ? ce08_mlX : 1'd0;
    assign ce14_mlB =
     invoke51_go_out ? ce09_mlX : 1'd0;
    assign ce14_reset = reset;
    assign ce15_addrA =
     invoke52_go_out ? ce010_addrX : 5'd0;
    assign ce15_addrB =
     invoke52_go_out ? ce011_addrX : 5'd0;
    assign ce15_clk = clk;
    assign ce15_go = invoke52_go_out;
    assign ce15_lenA =
     invoke52_go_out ? ce010_lenX : 5'd0;
    assign ce15_lenB =
     invoke52_go_out ? ce011_lenX : 5'd0;
    assign ce15_mlA =
     invoke52_go_out ? ce010_mlX : 1'd0;
    assign ce15_mlB =
     invoke52_go_out ? ce011_mlX : 1'd0;
    assign ce15_reset = reset;
    assign ce16_addrA =
     invoke53_go_out ? ce012_addrX : 5'd0;
    assign ce16_addrB =
     invoke53_go_out ? ce013_addrX : 5'd0;
    assign ce16_clk = clk;
    assign ce16_go = invoke53_go_out;
    assign ce16_lenA =
     invoke53_go_out ? ce012_lenX : 5'd0;
    assign ce16_lenB =
     invoke53_go_out ? ce013_lenX : 5'd0;
    assign ce16_mlA =
     invoke53_go_out ? ce012_mlX : 1'd0;
    assign ce16_mlB =
     invoke53_go_out ? ce013_mlX : 1'd0;
    assign ce16_reset = reset;
    assign ce17_addrA =
     invoke54_go_out ? ce014_addrX : 5'd0;
    assign ce17_addrB =
     invoke54_go_out ? ce015_addrX : 5'd0;
    assign ce17_clk = clk;
    assign ce17_go = invoke54_go_out;
    assign ce17_lenA =
     invoke54_go_out ? ce014_lenX : 5'd0;
    assign ce17_lenB =
     invoke54_go_out ? ce015_lenX : 5'd0;
    assign ce17_mlA =
     invoke54_go_out ? ce014_mlX : 1'd0;
    assign ce17_mlB =
     invoke54_go_out ? ce015_mlX : 1'd0;
    assign ce17_reset = reset;
    assign ce20_addrA =
     invoke55_go_out ? ce10_addrX : 5'd0;
    assign ce20_addrB =
     invoke55_go_out ? ce11_addrX : 5'd0;
    assign ce20_clk = clk;
    assign ce20_go = invoke55_go_out;
    assign ce20_lenA =
     invoke55_go_out ? ce10_lenX : 5'd0;
    assign ce20_lenB =
     invoke55_go_out ? ce11_lenX : 5'd0;
    assign ce20_mlA =
     invoke55_go_out ? ce10_mlX : 1'd0;
    assign ce20_mlB =
     invoke55_go_out ? ce11_mlX : 1'd0;
    assign ce20_reset = reset;
    assign ce21_addrA =
     invoke56_go_out ? ce12_addrX : 5'd0;
    assign ce21_addrB =
     invoke56_go_out ? ce13_addrX : 5'd0;
    assign ce21_clk = clk;
    assign ce21_go = invoke56_go_out;
    assign ce21_lenA =
     invoke56_go_out ? ce12_lenX : 5'd0;
    assign ce21_lenB =
     invoke56_go_out ? ce13_lenX : 5'd0;
    assign ce21_mlA =
     invoke56_go_out ? ce12_mlX : 1'd0;
    assign ce21_mlB =
     invoke56_go_out ? ce13_mlX : 1'd0;
    assign ce21_reset = reset;
    assign ce22_addrA =
     invoke57_go_out ? ce14_addrX : 5'd0;
    assign ce22_addrB =
     invoke57_go_out ? ce15_addrX : 5'd0;
    assign ce22_clk = clk;
    assign ce22_go = invoke57_go_out;
    assign ce22_lenA =
     invoke57_go_out ? ce14_lenX : 5'd0;
    assign ce22_lenB =
     invoke57_go_out ? ce15_lenX : 5'd0;
    assign ce22_mlA =
     invoke57_go_out ? ce14_mlX : 1'd0;
    assign ce22_mlB =
     invoke57_go_out ? ce15_mlX : 1'd0;
    assign ce22_reset = reset;
    assign ce23_addrA =
     invoke58_go_out ? ce16_addrX : 5'd0;
    assign ce23_addrB =
     invoke58_go_out ? ce17_addrX : 5'd0;
    assign ce23_clk = clk;
    assign ce23_go = invoke58_go_out;
    assign ce23_lenA =
     invoke58_go_out ? ce16_lenX : 5'd0;
    assign ce23_lenB =
     invoke58_go_out ? ce17_lenX : 5'd0;
    assign ce23_mlA =
     invoke58_go_out ? ce16_mlX : 1'd0;
    assign ce23_mlB =
     invoke58_go_out ? ce17_mlX : 1'd0;
    assign ce23_reset = reset;
    assign ce30_addrA =
     invoke59_go_out ? ce20_addrX : 5'd0;
    assign ce30_addrB =
     invoke59_go_out ? ce21_addrX : 5'd0;
    assign ce30_clk = clk;
    assign ce30_go = invoke59_go_out;
    assign ce30_lenA =
     invoke59_go_out ? ce20_lenX : 5'd0;
    assign ce30_lenB =
     invoke59_go_out ? ce21_lenX : 5'd0;
    assign ce30_mlA =
     invoke59_go_out ? ce20_mlX : 1'd0;
    assign ce30_mlB =
     invoke59_go_out ? ce21_mlX : 1'd0;
    assign ce30_reset = reset;
    assign ce31_addrA =
     invoke60_go_out ? ce22_addrX : 5'd0;
    assign ce31_addrB =
     invoke60_go_out ? ce23_addrX : 5'd0;
    assign ce31_clk = clk;
    assign ce31_go = invoke60_go_out;
    assign ce31_lenA =
     invoke60_go_out ? ce22_lenX : 5'd0;
    assign ce31_lenB =
     invoke60_go_out ? ce23_lenX : 5'd0;
    assign ce31_mlA =
     invoke60_go_out ? ce22_mlX : 1'd0;
    assign ce31_mlB =
     invoke60_go_out ? ce23_mlX : 1'd0;
    assign ce31_reset = reset;
    assign ce40_addrA =
     invoke61_go_out ? ce30_addrX : 5'd0;
    assign ce40_addrB =
     invoke61_go_out ? ce31_addrX : 5'd0;
    assign ce40_clk = clk;
    assign ce40_go = invoke61_go_out;
    assign ce40_lenA =
     invoke61_go_out ? ce30_lenX : 5'd0;
    assign ce40_lenB =
     invoke61_go_out ? ce31_lenX : 5'd0;
    assign ce40_mlA =
     invoke61_go_out ? ce30_mlX : 1'd0;
    assign ce40_mlB =
     invoke61_go_out ? ce31_mlX : 1'd0;
    assign ce40_reset = reset;
    assign comb_reg0_clk = clk;
    assign comb_reg0_in =
     find_write_index_go_out ? is_index0_out : 1'd0;
    assign comb_reg0_reset = reset;
    assign comb_reg0_write_en = find_write_index_go_out;
    assign comb_reg1_clk = clk;
    assign comb_reg1_in =
     find_write_index_go_out ? is_index1_out :
     is_length_zero0_go_out ? z_eq_out : 1'd0;
    assign comb_reg1_reset = reset;
    assign comb_reg1_write_en = find_write_index_go_out | is_length_zero0_go_out;
    assign comb_reg10_clk = clk;
    assign comb_reg10_in =
     find_write_index_go_out ? is_index10_out : 1'd0;
    assign comb_reg10_reset = reset;
    assign comb_reg10_write_en = find_write_index_go_out;
    assign comb_reg11_clk = clk;
    assign comb_reg11_in =
     find_write_index_go_out ? is_index11_out : 1'd0;
    assign comb_reg11_reset = reset;
    assign comb_reg11_write_en = find_write_index_go_out;
    assign comb_reg12_clk = clk;
    assign comb_reg12_in =
     find_write_index_go_out ? is_index12_out : 1'd0;
    assign comb_reg12_reset = reset;
    assign comb_reg12_write_en = find_write_index_go_out;
    assign comb_reg13_clk = clk;
    assign comb_reg13_in =
     find_write_index_go_out ? is_index13_out : 1'd0;
    assign comb_reg13_reset = reset;
    assign comb_reg13_write_en = find_write_index_go_out;
    assign comb_reg14_clk = clk;
    assign comb_reg14_in =
     find_write_index_go_out ? is_index14_out : 1'd0;
    assign comb_reg14_reset = reset;
    assign comb_reg14_write_en = find_write_index_go_out;
    assign comb_reg15_clk = clk;
    assign comb_reg15_in =
     find_write_index_go_out ? is_index15_out : 1'd0;
    assign comb_reg15_reset = reset;
    assign comb_reg15_write_en = find_write_index_go_out;
    assign comb_reg16_clk = clk;
    assign comb_reg16_in =
     find_write_index_go_out ? is_index16_out : 1'd0;
    assign comb_reg16_reset = reset;
    assign comb_reg16_write_en = find_write_index_go_out;
    assign comb_reg17_clk = clk;
    assign comb_reg17_in =
     find_write_index_go_out ? is_index17_out : 1'd0;
    assign comb_reg17_reset = reset;
    assign comb_reg17_write_en = find_write_index_go_out;
    assign comb_reg18_clk = clk;
    assign comb_reg18_in =
     find_write_index_go_out ? is_index18_out : 1'd0;
    assign comb_reg18_reset = reset;
    assign comb_reg18_write_en = find_write_index_go_out;
    assign comb_reg19_clk = clk;
    assign comb_reg19_in =
     find_write_index_go_out ? is_index19_out : 1'd0;
    assign comb_reg19_reset = reset;
    assign comb_reg19_write_en = find_write_index_go_out;
    assign comb_reg2_clk = clk;
    assign comb_reg2_in =
     find_write_index_go_out ? is_index2_out : 1'd0;
    assign comb_reg2_reset = reset;
    assign comb_reg2_write_en = find_write_index_go_out;
    assign comb_reg20_clk = clk;
    assign comb_reg20_in =
     find_write_index_go_out ? is_index20_out : 1'd0;
    assign comb_reg20_reset = reset;
    assign comb_reg20_write_en = find_write_index_go_out;
    assign comb_reg21_clk = clk;
    assign comb_reg21_in =
     find_write_index_go_out ? is_index21_out : 1'd0;
    assign comb_reg21_reset = reset;
    assign comb_reg21_write_en = find_write_index_go_out;
    assign comb_reg22_clk = clk;
    assign comb_reg22_in =
     find_write_index_go_out ? is_index22_out : 1'd0;
    assign comb_reg22_reset = reset;
    assign comb_reg22_write_en = find_write_index_go_out;
    assign comb_reg23_clk = clk;
    assign comb_reg23_in =
     find_write_index_go_out ? is_index23_out : 1'd0;
    assign comb_reg23_reset = reset;
    assign comb_reg23_write_en = find_write_index_go_out;
    assign comb_reg24_clk = clk;
    assign comb_reg24_in =
     find_write_index_go_out ? is_index24_out : 1'd0;
    assign comb_reg24_reset = reset;
    assign comb_reg24_write_en = find_write_index_go_out;
    assign comb_reg25_clk = clk;
    assign comb_reg25_in =
     find_write_index_go_out ? is_index25_out : 1'd0;
    assign comb_reg25_reset = reset;
    assign comb_reg25_write_en = find_write_index_go_out;
    assign comb_reg26_clk = clk;
    assign comb_reg26_in =
     find_write_index_go_out ? is_index26_out : 1'd0;
    assign comb_reg26_reset = reset;
    assign comb_reg26_write_en = find_write_index_go_out;
    assign comb_reg27_clk = clk;
    assign comb_reg27_in =
     find_write_index_go_out ? is_index27_out : 1'd0;
    assign comb_reg27_reset = reset;
    assign comb_reg27_write_en = find_write_index_go_out;
    assign comb_reg28_clk = clk;
    assign comb_reg28_in =
     find_write_index_go_out ? is_index28_out : 1'd0;
    assign comb_reg28_reset = reset;
    assign comb_reg28_write_en = find_write_index_go_out;
    assign comb_reg29_clk = clk;
    assign comb_reg29_in =
     find_write_index_go_out ? is_index29_out : 1'd0;
    assign comb_reg29_reset = reset;
    assign comb_reg29_write_en = find_write_index_go_out;
    assign comb_reg3_clk = clk;
    assign comb_reg3_in =
     find_write_index_go_out ? is_index3_out : 1'd0;
    assign comb_reg3_reset = reset;
    assign comb_reg3_write_en = find_write_index_go_out;
    assign comb_reg30_clk = clk;
    assign comb_reg30_in =
     find_write_index_go_out ? is_index30_out : 1'd0;
    assign comb_reg30_reset = reset;
    assign comb_reg30_write_en = find_write_index_go_out;
    assign comb_reg31_clk = clk;
    assign comb_reg31_in =
     find_write_index_go_out ? is_index31_out : 1'd0;
    assign comb_reg31_reset = reset;
    assign comb_reg31_write_en = find_write_index_go_out;
    assign comb_reg4_clk = clk;
    assign comb_reg4_in =
     find_write_index_go_out ? is_index4_out : 1'd0;
    assign comb_reg4_reset = reset;
    assign comb_reg4_write_en = find_write_index_go_out;
    assign comb_reg5_clk = clk;
    assign comb_reg5_in =
     find_write_index_go_out ? is_index5_out : 1'd0;
    assign comb_reg5_reset = reset;
    assign comb_reg5_write_en = find_write_index_go_out;
    assign comb_reg6_clk = clk;
    assign comb_reg6_in =
     find_write_index_go_out ? is_index6_out : 1'd0;
    assign comb_reg6_reset = reset;
    assign comb_reg6_write_en = find_write_index_go_out;
    assign comb_reg7_clk = clk;
    assign comb_reg7_in =
     find_write_index_go_out ? is_index7_out : 1'd0;
    assign comb_reg7_reset = reset;
    assign comb_reg7_write_en = find_write_index_go_out;
    assign comb_reg8_clk = clk;
    assign comb_reg8_in =
     find_write_index_go_out ? is_index8_out : 1'd0;
    assign comb_reg8_reset = reset;
    assign comb_reg8_write_en = find_write_index_go_out;
    assign comb_reg9_clk = clk;
    assign comb_reg9_in =
     find_write_index_go_out ? is_index9_out : 1'd0;
    assign comb_reg9_reset = reset;
    assign comb_reg9_write_en = find_write_index_go_out;
    assign default_to_zero_length_index_done_in = out_done;
    assign default_to_zero_length_index_go_in = ~default_to_zero_length_index_done_out & fsm32_out == 4'd8 & tdcc32_go_out;
    assign find_write_index_done_in = comb_reg0_done;
    assign find_write_index_go_in = ~find_write_index_done_out & fsm31_out == 3'd3 & tdcc31_go_out;
    assign fsm_clk = clk;
    assign fsm_in =
     fsm_out == 2'd2 ? 2'd0 :
     fsm_out == 2'd0 & comb_reg0_out & tdcc_go_out ? 2'd1 :
     fsm_out == 2'd1 & write0_done_out & tdcc_go_out | fsm_out == 2'd0 & ~comb_reg0_out & tdcc_go_out ? 2'd2 : 2'd0;
    assign fsm_reset = reset;
    assign fsm_write_en = fsm_out == 2'd2 | fsm_out == 2'd0 & comb_reg0_out & tdcc_go_out | fsm_out == 2'd1 & write0_done_out & tdcc_go_out | fsm_out == 2'd0 & ~comb_reg0_out & tdcc_go_out;
    assign fsm0_clk = clk;
    assign fsm0_in =
     fsm0_out == 2'd2 ? 2'd0 :
     fsm0_out == 2'd0 & comb_reg1_out & tdcc0_go_out ? 2'd1 :
     fsm0_out == 2'd1 & write1_done_out & tdcc0_go_out | fsm0_out == 2'd0 & ~comb_reg1_out & tdcc0_go_out ? 2'd2 : 2'd0;
    assign fsm0_reset = reset;
    assign fsm0_write_en = fsm0_out == 2'd2 | fsm0_out == 2'd0 & comb_reg1_out & tdcc0_go_out | fsm0_out == 2'd1 & write1_done_out & tdcc0_go_out | fsm0_out == 2'd0 & ~comb_reg1_out & tdcc0_go_out;
    assign fsm1_clk = clk;
    assign fsm1_in =
     fsm1_out == 2'd2 ? 2'd0 :
     fsm1_out == 2'd0 & comb_reg2_out & tdcc1_go_out ? 2'd1 :
     fsm1_out == 2'd1 & write2_done_out & tdcc1_go_out | fsm1_out == 2'd0 & ~comb_reg2_out & tdcc1_go_out ? 2'd2 : 2'd0;
    assign fsm1_reset = reset;
    assign fsm1_write_en = fsm1_out == 2'd2 | fsm1_out == 2'd0 & comb_reg2_out & tdcc1_go_out | fsm1_out == 2'd1 & write2_done_out & tdcc1_go_out | fsm1_out == 2'd0 & ~comb_reg2_out & tdcc1_go_out;
    assign fsm10_clk = clk;
    assign fsm10_in =
     fsm10_out == 2'd2 ? 2'd0 :
     fsm10_out == 2'd0 & comb_reg11_out & tdcc10_go_out ? 2'd1 :
     fsm10_out == 2'd1 & write11_done_out & tdcc10_go_out | fsm10_out == 2'd0 & ~comb_reg11_out & tdcc10_go_out ? 2'd2 : 2'd0;
    assign fsm10_reset = reset;
    assign fsm10_write_en = fsm10_out == 2'd2 | fsm10_out == 2'd0 & comb_reg11_out & tdcc10_go_out | fsm10_out == 2'd1 & write11_done_out & tdcc10_go_out | fsm10_out == 2'd0 & ~comb_reg11_out & tdcc10_go_out;
    assign fsm11_clk = clk;
    assign fsm11_in =
     fsm11_out == 2'd2 ? 2'd0 :
     fsm11_out == 2'd0 & comb_reg12_out & tdcc11_go_out ? 2'd1 :
     fsm11_out == 2'd1 & write12_done_out & tdcc11_go_out | fsm11_out == 2'd0 & ~comb_reg12_out & tdcc11_go_out ? 2'd2 : 2'd0;
    assign fsm11_reset = reset;
    assign fsm11_write_en = fsm11_out == 2'd2 | fsm11_out == 2'd0 & comb_reg12_out & tdcc11_go_out | fsm11_out == 2'd1 & write12_done_out & tdcc11_go_out | fsm11_out == 2'd0 & ~comb_reg12_out & tdcc11_go_out;
    assign fsm12_clk = clk;
    assign fsm12_in =
     fsm12_out == 2'd2 ? 2'd0 :
     fsm12_out == 2'd0 & comb_reg13_out & tdcc12_go_out ? 2'd1 :
     fsm12_out == 2'd1 & write13_done_out & tdcc12_go_out | fsm12_out == 2'd0 & ~comb_reg13_out & tdcc12_go_out ? 2'd2 : 2'd0;
    assign fsm12_reset = reset;
    assign fsm12_write_en = fsm12_out == 2'd2 | fsm12_out == 2'd0 & comb_reg13_out & tdcc12_go_out | fsm12_out == 2'd1 & write13_done_out & tdcc12_go_out | fsm12_out == 2'd0 & ~comb_reg13_out & tdcc12_go_out;
    assign fsm13_clk = clk;
    assign fsm13_in =
     fsm13_out == 2'd2 ? 2'd0 :
     fsm13_out == 2'd0 & comb_reg14_out & tdcc13_go_out ? 2'd1 :
     fsm13_out == 2'd1 & write14_done_out & tdcc13_go_out | fsm13_out == 2'd0 & ~comb_reg14_out & tdcc13_go_out ? 2'd2 : 2'd0;
    assign fsm13_reset = reset;
    assign fsm13_write_en = fsm13_out == 2'd2 | fsm13_out == 2'd0 & comb_reg14_out & tdcc13_go_out | fsm13_out == 2'd1 & write14_done_out & tdcc13_go_out | fsm13_out == 2'd0 & ~comb_reg14_out & tdcc13_go_out;
    assign fsm14_clk = clk;
    assign fsm14_in =
     fsm14_out == 2'd2 ? 2'd0 :
     fsm14_out == 2'd0 & comb_reg15_out & tdcc14_go_out ? 2'd1 :
     fsm14_out == 2'd1 & write15_done_out & tdcc14_go_out | fsm14_out == 2'd0 & ~comb_reg15_out & tdcc14_go_out ? 2'd2 : 2'd0;
    assign fsm14_reset = reset;
    assign fsm14_write_en = fsm14_out == 2'd2 | fsm14_out == 2'd0 & comb_reg15_out & tdcc14_go_out | fsm14_out == 2'd1 & write15_done_out & tdcc14_go_out | fsm14_out == 2'd0 & ~comb_reg15_out & tdcc14_go_out;
    assign fsm15_clk = clk;
    assign fsm15_in =
     fsm15_out == 2'd2 ? 2'd0 :
     fsm15_out == 2'd0 & comb_reg16_out & tdcc15_go_out ? 2'd1 :
     fsm15_out == 2'd1 & write16_done_out & tdcc15_go_out | fsm15_out == 2'd0 & ~comb_reg16_out & tdcc15_go_out ? 2'd2 : 2'd0;
    assign fsm15_reset = reset;
    assign fsm15_write_en = fsm15_out == 2'd2 | fsm15_out == 2'd0 & comb_reg16_out & tdcc15_go_out | fsm15_out == 2'd1 & write16_done_out & tdcc15_go_out | fsm15_out == 2'd0 & ~comb_reg16_out & tdcc15_go_out;
    assign fsm16_clk = clk;
    assign fsm16_in =
     fsm16_out == 2'd2 ? 2'd0 :
     fsm16_out == 2'd0 & comb_reg17_out & tdcc16_go_out ? 2'd1 :
     fsm16_out == 2'd1 & write17_done_out & tdcc16_go_out | fsm16_out == 2'd0 & ~comb_reg17_out & tdcc16_go_out ? 2'd2 : 2'd0;
    assign fsm16_reset = reset;
    assign fsm16_write_en = fsm16_out == 2'd2 | fsm16_out == 2'd0 & comb_reg17_out & tdcc16_go_out | fsm16_out == 2'd1 & write17_done_out & tdcc16_go_out | fsm16_out == 2'd0 & ~comb_reg17_out & tdcc16_go_out;
    assign fsm17_clk = clk;
    assign fsm17_in =
     fsm17_out == 2'd2 ? 2'd0 :
     fsm17_out == 2'd0 & comb_reg18_out & tdcc17_go_out ? 2'd1 :
     fsm17_out == 2'd1 & write18_done_out & tdcc17_go_out | fsm17_out == 2'd0 & ~comb_reg18_out & tdcc17_go_out ? 2'd2 : 2'd0;
    assign fsm17_reset = reset;
    assign fsm17_write_en = fsm17_out == 2'd2 | fsm17_out == 2'd0 & comb_reg18_out & tdcc17_go_out | fsm17_out == 2'd1 & write18_done_out & tdcc17_go_out | fsm17_out == 2'd0 & ~comb_reg18_out & tdcc17_go_out;
    assign fsm18_clk = clk;
    assign fsm18_in =
     fsm18_out == 2'd2 ? 2'd0 :
     fsm18_out == 2'd0 & comb_reg19_out & tdcc18_go_out ? 2'd1 :
     fsm18_out == 2'd1 & write19_done_out & tdcc18_go_out | fsm18_out == 2'd0 & ~comb_reg19_out & tdcc18_go_out ? 2'd2 : 2'd0;
    assign fsm18_reset = reset;
    assign fsm18_write_en = fsm18_out == 2'd2 | fsm18_out == 2'd0 & comb_reg19_out & tdcc18_go_out | fsm18_out == 2'd1 & write19_done_out & tdcc18_go_out | fsm18_out == 2'd0 & ~comb_reg19_out & tdcc18_go_out;
    assign fsm19_clk = clk;
    assign fsm19_in =
     fsm19_out == 2'd2 ? 2'd0 :
     fsm19_out == 2'd0 & comb_reg20_out & tdcc19_go_out ? 2'd1 :
     fsm19_out == 2'd1 & write20_done_out & tdcc19_go_out | fsm19_out == 2'd0 & ~comb_reg20_out & tdcc19_go_out ? 2'd2 : 2'd0;
    assign fsm19_reset = reset;
    assign fsm19_write_en = fsm19_out == 2'd2 | fsm19_out == 2'd0 & comb_reg20_out & tdcc19_go_out | fsm19_out == 2'd1 & write20_done_out & tdcc19_go_out | fsm19_out == 2'd0 & ~comb_reg20_out & tdcc19_go_out;
    assign fsm2_clk = clk;
    assign fsm2_in =
     fsm2_out == 2'd2 ? 2'd0 :
     fsm2_out == 2'd0 & comb_reg3_out & tdcc2_go_out ? 2'd1 :
     fsm2_out == 2'd1 & write3_done_out & tdcc2_go_out | fsm2_out == 2'd0 & ~comb_reg3_out & tdcc2_go_out ? 2'd2 : 2'd0;
    assign fsm2_reset = reset;
    assign fsm2_write_en = fsm2_out == 2'd2 | fsm2_out == 2'd0 & comb_reg3_out & tdcc2_go_out | fsm2_out == 2'd1 & write3_done_out & tdcc2_go_out | fsm2_out == 2'd0 & ~comb_reg3_out & tdcc2_go_out;
    assign fsm20_clk = clk;
    assign fsm20_in =
     fsm20_out == 2'd2 ? 2'd0 :
     fsm20_out == 2'd0 & comb_reg21_out & tdcc20_go_out ? 2'd1 :
     fsm20_out == 2'd1 & write21_done_out & tdcc20_go_out | fsm20_out == 2'd0 & ~comb_reg21_out & tdcc20_go_out ? 2'd2 : 2'd0;
    assign fsm20_reset = reset;
    assign fsm20_write_en = fsm20_out == 2'd2 | fsm20_out == 2'd0 & comb_reg21_out & tdcc20_go_out | fsm20_out == 2'd1 & write21_done_out & tdcc20_go_out | fsm20_out == 2'd0 & ~comb_reg21_out & tdcc20_go_out;
    assign fsm21_clk = clk;
    assign fsm21_in =
     fsm21_out == 2'd2 ? 2'd0 :
     fsm21_out == 2'd0 & comb_reg22_out & tdcc21_go_out ? 2'd1 :
     fsm21_out == 2'd1 & write22_done_out & tdcc21_go_out | fsm21_out == 2'd0 & ~comb_reg22_out & tdcc21_go_out ? 2'd2 : 2'd0;
    assign fsm21_reset = reset;
    assign fsm21_write_en = fsm21_out == 2'd2 | fsm21_out == 2'd0 & comb_reg22_out & tdcc21_go_out | fsm21_out == 2'd1 & write22_done_out & tdcc21_go_out | fsm21_out == 2'd0 & ~comb_reg22_out & tdcc21_go_out;
    assign fsm22_clk = clk;
    assign fsm22_in =
     fsm22_out == 2'd2 ? 2'd0 :
     fsm22_out == 2'd0 & comb_reg23_out & tdcc22_go_out ? 2'd1 :
     fsm22_out == 2'd1 & write23_done_out & tdcc22_go_out | fsm22_out == 2'd0 & ~comb_reg23_out & tdcc22_go_out ? 2'd2 : 2'd0;
    assign fsm22_reset = reset;
    assign fsm22_write_en = fsm22_out == 2'd2 | fsm22_out == 2'd0 & comb_reg23_out & tdcc22_go_out | fsm22_out == 2'd1 & write23_done_out & tdcc22_go_out | fsm22_out == 2'd0 & ~comb_reg23_out & tdcc22_go_out;
    assign fsm23_clk = clk;
    assign fsm23_in =
     fsm23_out == 2'd2 ? 2'd0 :
     fsm23_out == 2'd0 & comb_reg24_out & tdcc23_go_out ? 2'd1 :
     fsm23_out == 2'd1 & write24_done_out & tdcc23_go_out | fsm23_out == 2'd0 & ~comb_reg24_out & tdcc23_go_out ? 2'd2 : 2'd0;
    assign fsm23_reset = reset;
    assign fsm23_write_en = fsm23_out == 2'd2 | fsm23_out == 2'd0 & comb_reg24_out & tdcc23_go_out | fsm23_out == 2'd1 & write24_done_out & tdcc23_go_out | fsm23_out == 2'd0 & ~comb_reg24_out & tdcc23_go_out;
    assign fsm24_clk = clk;
    assign fsm24_in =
     fsm24_out == 2'd2 ? 2'd0 :
     fsm24_out == 2'd0 & comb_reg25_out & tdcc24_go_out ? 2'd1 :
     fsm24_out == 2'd1 & write25_done_out & tdcc24_go_out | fsm24_out == 2'd0 & ~comb_reg25_out & tdcc24_go_out ? 2'd2 : 2'd0;
    assign fsm24_reset = reset;
    assign fsm24_write_en = fsm24_out == 2'd2 | fsm24_out == 2'd0 & comb_reg25_out & tdcc24_go_out | fsm24_out == 2'd1 & write25_done_out & tdcc24_go_out | fsm24_out == 2'd0 & ~comb_reg25_out & tdcc24_go_out;
    assign fsm25_clk = clk;
    assign fsm25_in =
     fsm25_out == 2'd2 ? 2'd0 :
     fsm25_out == 2'd0 & comb_reg26_out & tdcc25_go_out ? 2'd1 :
     fsm25_out == 2'd1 & write26_done_out & tdcc25_go_out | fsm25_out == 2'd0 & ~comb_reg26_out & tdcc25_go_out ? 2'd2 : 2'd0;
    assign fsm25_reset = reset;
    assign fsm25_write_en = fsm25_out == 2'd2 | fsm25_out == 2'd0 & comb_reg26_out & tdcc25_go_out | fsm25_out == 2'd1 & write26_done_out & tdcc25_go_out | fsm25_out == 2'd0 & ~comb_reg26_out & tdcc25_go_out;
    assign fsm26_clk = clk;
    assign fsm26_in =
     fsm26_out == 2'd2 ? 2'd0 :
     fsm26_out == 2'd0 & comb_reg27_out & tdcc26_go_out ? 2'd1 :
     fsm26_out == 2'd1 & write27_done_out & tdcc26_go_out | fsm26_out == 2'd0 & ~comb_reg27_out & tdcc26_go_out ? 2'd2 : 2'd0;
    assign fsm26_reset = reset;
    assign fsm26_write_en = fsm26_out == 2'd2 | fsm26_out == 2'd0 & comb_reg27_out & tdcc26_go_out | fsm26_out == 2'd1 & write27_done_out & tdcc26_go_out | fsm26_out == 2'd0 & ~comb_reg27_out & tdcc26_go_out;
    assign fsm27_clk = clk;
    assign fsm27_in =
     fsm27_out == 2'd2 ? 2'd0 :
     fsm27_out == 2'd0 & comb_reg28_out & tdcc27_go_out ? 2'd1 :
     fsm27_out == 2'd1 & write28_done_out & tdcc27_go_out | fsm27_out == 2'd0 & ~comb_reg28_out & tdcc27_go_out ? 2'd2 : 2'd0;
    assign fsm27_reset = reset;
    assign fsm27_write_en = fsm27_out == 2'd2 | fsm27_out == 2'd0 & comb_reg28_out & tdcc27_go_out | fsm27_out == 2'd1 & write28_done_out & tdcc27_go_out | fsm27_out == 2'd0 & ~comb_reg28_out & tdcc27_go_out;
    assign fsm28_clk = clk;
    assign fsm28_in =
     fsm28_out == 2'd2 ? 2'd0 :
     fsm28_out == 2'd0 & comb_reg29_out & tdcc28_go_out ? 2'd1 :
     fsm28_out == 2'd1 & write29_done_out & tdcc28_go_out | fsm28_out == 2'd0 & ~comb_reg29_out & tdcc28_go_out ? 2'd2 : 2'd0;
    assign fsm28_reset = reset;
    assign fsm28_write_en = fsm28_out == 2'd2 | fsm28_out == 2'd0 & comb_reg29_out & tdcc28_go_out | fsm28_out == 2'd1 & write29_done_out & tdcc28_go_out | fsm28_out == 2'd0 & ~comb_reg29_out & tdcc28_go_out;
    assign fsm29_clk = clk;
    assign fsm29_in =
     fsm29_out == 2'd2 ? 2'd0 :
     fsm29_out == 2'd0 & comb_reg30_out & tdcc29_go_out ? 2'd1 :
     fsm29_out == 2'd1 & write30_done_out & tdcc29_go_out | fsm29_out == 2'd0 & ~comb_reg30_out & tdcc29_go_out ? 2'd2 : 2'd0;
    assign fsm29_reset = reset;
    assign fsm29_write_en = fsm29_out == 2'd2 | fsm29_out == 2'd0 & comb_reg30_out & tdcc29_go_out | fsm29_out == 2'd1 & write30_done_out & tdcc29_go_out | fsm29_out == 2'd0 & ~comb_reg30_out & tdcc29_go_out;
    assign fsm3_clk = clk;
    assign fsm3_in =
     fsm3_out == 2'd2 ? 2'd0 :
     fsm3_out == 2'd0 & comb_reg4_out & tdcc3_go_out ? 2'd1 :
     fsm3_out == 2'd1 & write4_done_out & tdcc3_go_out | fsm3_out == 2'd0 & ~comb_reg4_out & tdcc3_go_out ? 2'd2 : 2'd0;
    assign fsm3_reset = reset;
    assign fsm3_write_en = fsm3_out == 2'd2 | fsm3_out == 2'd0 & comb_reg4_out & tdcc3_go_out | fsm3_out == 2'd1 & write4_done_out & tdcc3_go_out | fsm3_out == 2'd0 & ~comb_reg4_out & tdcc3_go_out;
    assign fsm30_clk = clk;
    assign fsm30_in =
     fsm30_out == 2'd2 ? 2'd0 :
     fsm30_out == 2'd0 & comb_reg31_out & tdcc30_go_out ? 2'd1 :
     fsm30_out == 2'd1 & write31_done_out & tdcc30_go_out | fsm30_out == 2'd0 & ~comb_reg31_out & tdcc30_go_out ? 2'd2 : 2'd0;
    assign fsm30_reset = reset;
    assign fsm30_write_en = fsm30_out == 2'd2 | fsm30_out == 2'd0 & comb_reg31_out & tdcc30_go_out | fsm30_out == 2'd1 & write31_done_out & tdcc30_go_out | fsm30_out == 2'd0 & ~comb_reg31_out & tdcc30_go_out;
    assign fsm31_clk = clk;
    assign fsm31_in =
     fsm31_out == 3'd5 ? 3'd0 :
     fsm31_out == 3'd0 & write_en & tdcc31_go_out ? 3'd1 :
     fsm31_out == 3'd1 & is_length_zero0_done_out & comb_reg1_out & tdcc31_go_out ? 3'd2 :
     fsm31_out == 3'd1 & is_length_zero0_done_out & ~comb_reg1_out & tdcc31_go_out ? 3'd3 :
     fsm31_out == 3'd3 & find_write_index_done_out & tdcc31_go_out ? 3'd4 :
     fsm31_out == 3'd2 & write_zero_done_out & tdcc31_go_out | fsm31_out == 3'd4 & par_done_out & tdcc31_go_out | fsm31_out == 3'd0 & ~write_en & tdcc31_go_out ? 3'd5 : 3'd0;
    assign fsm31_reset = reset;
    assign fsm31_write_en = fsm31_out == 3'd5 | fsm31_out == 3'd0 & write_en & tdcc31_go_out | fsm31_out == 3'd1 & is_length_zero0_done_out & comb_reg1_out & tdcc31_go_out | fsm31_out == 3'd1 & is_length_zero0_done_out & ~comb_reg1_out & tdcc31_go_out | fsm31_out == 3'd3 & find_write_index_done_out & tdcc31_go_out | fsm31_out == 3'd2 & write_zero_done_out & tdcc31_go_out | fsm31_out == 3'd4 & par_done_out & tdcc31_go_out | fsm31_out == 3'd0 & ~write_en & tdcc31_go_out;
    assign fsm32_clk = clk;
    assign fsm32_in =
     fsm32_out == 4'd9 ? 4'd0 :
     fsm32_out == 4'd0 & search_en & tdcc32_go_out ? 4'd1 :
     fsm32_out == 4'd1 & par0_done_out & tdcc32_go_out ? 4'd2 :
     fsm32_out == 4'd2 & par1_done_out & tdcc32_go_out ? 4'd3 :
     fsm32_out == 4'd3 & par2_done_out & tdcc32_go_out ? 4'd4 :
     fsm32_out == 4'd4 & par3_done_out & tdcc32_go_out ? 4'd5 :
     fsm32_out == 4'd5 & par4_done_out & tdcc32_go_out ? 4'd6 :
     fsm32_out == 4'd6 & invoke61_done_out & ce40_mlX & tdcc32_go_out ? 4'd7 :
     fsm32_out == 4'd6 & invoke61_done_out & ~ce40_mlX & tdcc32_go_out ? 4'd8 :
     fsm32_out == 4'd7 & save_index_done_out & tdcc32_go_out | fsm32_out == 4'd8 & default_to_zero_length_index_done_out & tdcc32_go_out | fsm32_out == 4'd0 & ~search_en & tdcc32_go_out ? 4'd9 : 4'd0;
    assign fsm32_reset = reset;
    assign fsm32_write_en = fsm32_out == 4'd9 | fsm32_out == 4'd0 & search_en & tdcc32_go_out | fsm32_out == 4'd1 & par0_done_out & tdcc32_go_out | fsm32_out == 4'd2 & par1_done_out & tdcc32_go_out | fsm32_out == 4'd3 & par2_done_out & tdcc32_go_out | fsm32_out == 4'd4 & par3_done_out & tdcc32_go_out | fsm32_out == 4'd5 & par4_done_out & tdcc32_go_out | fsm32_out == 4'd6 & invoke61_done_out & ce40_mlX & tdcc32_go_out | fsm32_out == 4'd6 & invoke61_done_out & ~ce40_mlX & tdcc32_go_out | fsm32_out == 4'd7 & save_index_done_out & tdcc32_go_out | fsm32_out == 4'd8 & default_to_zero_length_index_done_out & tdcc32_go_out | fsm32_out == 4'd0 & ~search_en & tdcc32_go_out;
    assign fsm33_clk = clk;
    assign fsm33_in =
     fsm33_out == 1'd1 ? 1'd0 :
     fsm33_out == 1'd0 & par5_done_out & tdcc33_go_out ? 1'd1 : 1'd0;
    assign fsm33_reset = reset;
    assign fsm33_write_en = fsm33_out == 1'd1 | fsm33_out == 1'd0 & par5_done_out & tdcc33_go_out;
    assign fsm4_clk = clk;
    assign fsm4_in =
     fsm4_out == 2'd2 ? 2'd0 :
     fsm4_out == 2'd0 & comb_reg5_out & tdcc4_go_out ? 2'd1 :
     fsm4_out == 2'd1 & write5_done_out & tdcc4_go_out | fsm4_out == 2'd0 & ~comb_reg5_out & tdcc4_go_out ? 2'd2 : 2'd0;
    assign fsm4_reset = reset;
    assign fsm4_write_en = fsm4_out == 2'd2 | fsm4_out == 2'd0 & comb_reg5_out & tdcc4_go_out | fsm4_out == 2'd1 & write5_done_out & tdcc4_go_out | fsm4_out == 2'd0 & ~comb_reg5_out & tdcc4_go_out;
    assign fsm5_clk = clk;
    assign fsm5_in =
     fsm5_out == 2'd2 ? 2'd0 :
     fsm5_out == 2'd0 & comb_reg6_out & tdcc5_go_out ? 2'd1 :
     fsm5_out == 2'd1 & write6_done_out & tdcc5_go_out | fsm5_out == 2'd0 & ~comb_reg6_out & tdcc5_go_out ? 2'd2 : 2'd0;
    assign fsm5_reset = reset;
    assign fsm5_write_en = fsm5_out == 2'd2 | fsm5_out == 2'd0 & comb_reg6_out & tdcc5_go_out | fsm5_out == 2'd1 & write6_done_out & tdcc5_go_out | fsm5_out == 2'd0 & ~comb_reg6_out & tdcc5_go_out;
    assign fsm6_clk = clk;
    assign fsm6_in =
     fsm6_out == 2'd2 ? 2'd0 :
     fsm6_out == 2'd0 & comb_reg7_out & tdcc6_go_out ? 2'd1 :
     fsm6_out == 2'd1 & write7_done_out & tdcc6_go_out | fsm6_out == 2'd0 & ~comb_reg7_out & tdcc6_go_out ? 2'd2 : 2'd0;
    assign fsm6_reset = reset;
    assign fsm6_write_en = fsm6_out == 2'd2 | fsm6_out == 2'd0 & comb_reg7_out & tdcc6_go_out | fsm6_out == 2'd1 & write7_done_out & tdcc6_go_out | fsm6_out == 2'd0 & ~comb_reg7_out & tdcc6_go_out;
    assign fsm7_clk = clk;
    assign fsm7_in =
     fsm7_out == 2'd2 ? 2'd0 :
     fsm7_out == 2'd0 & comb_reg8_out & tdcc7_go_out ? 2'd1 :
     fsm7_out == 2'd1 & write8_done_out & tdcc7_go_out | fsm7_out == 2'd0 & ~comb_reg8_out & tdcc7_go_out ? 2'd2 : 2'd0;
    assign fsm7_reset = reset;
    assign fsm7_write_en = fsm7_out == 2'd2 | fsm7_out == 2'd0 & comb_reg8_out & tdcc7_go_out | fsm7_out == 2'd1 & write8_done_out & tdcc7_go_out | fsm7_out == 2'd0 & ~comb_reg8_out & tdcc7_go_out;
    assign fsm8_clk = clk;
    assign fsm8_in =
     fsm8_out == 2'd2 ? 2'd0 :
     fsm8_out == 2'd0 & comb_reg9_out & tdcc8_go_out ? 2'd1 :
     fsm8_out == 2'd1 & write9_done_out & tdcc8_go_out | fsm8_out == 2'd0 & ~comb_reg9_out & tdcc8_go_out ? 2'd2 : 2'd0;
    assign fsm8_reset = reset;
    assign fsm8_write_en = fsm8_out == 2'd2 | fsm8_out == 2'd0 & comb_reg9_out & tdcc8_go_out | fsm8_out == 2'd1 & write9_done_out & tdcc8_go_out | fsm8_out == 2'd0 & ~comb_reg9_out & tdcc8_go_out;
    assign fsm9_clk = clk;
    assign fsm9_in =
     fsm9_out == 2'd2 ? 2'd0 :
     fsm9_out == 2'd0 & comb_reg10_out & tdcc9_go_out ? 2'd1 :
     fsm9_out == 2'd1 & write10_done_out & tdcc9_go_out | fsm9_out == 2'd0 & ~comb_reg10_out & tdcc9_go_out ? 2'd2 : 2'd0;
    assign fsm9_reset = reset;
    assign fsm9_write_en = fsm9_out == 2'd2 | fsm9_out == 2'd0 & comb_reg10_out & tdcc9_go_out | fsm9_out == 2'd1 & write10_done_out & tdcc9_go_out | fsm9_out == 2'd0 & ~comb_reg10_out & tdcc9_go_out;
    assign invoke0_done_in = me1_done;
    assign invoke0_go_in = ~(pd32_out | invoke0_done_out) & par0_go_out;
    assign invoke10_done_in = me11_done;
    assign invoke10_go_in = ~(pd42_out | invoke10_done_out) & par0_go_out;
    assign invoke11_done_in = me12_done;
    assign invoke11_go_in = ~(pd43_out | invoke11_done_out) & par0_go_out;
    assign invoke12_done_in = me13_done;
    assign invoke12_go_in = ~(pd44_out | invoke12_done_out) & par0_go_out;
    assign invoke13_done_in = me14_done;
    assign invoke13_go_in = ~(pd45_out | invoke13_done_out) & par0_go_out;
    assign invoke14_done_in = me15_done;
    assign invoke14_go_in = ~(pd46_out | invoke14_done_out) & par0_go_out;
    assign invoke15_done_in = me16_done;
    assign invoke15_go_in = ~(pd47_out | invoke15_done_out) & par0_go_out;
    assign invoke16_done_in = me17_done;
    assign invoke16_go_in = ~(pd48_out | invoke16_done_out) & par0_go_out;
    assign invoke17_done_in = me18_done;
    assign invoke17_go_in = ~(pd49_out | invoke17_done_out) & par0_go_out;
    assign invoke18_done_in = me19_done;
    assign invoke18_go_in = ~(pd50_out | invoke18_done_out) & par0_go_out;
    assign invoke19_done_in = me20_done;
    assign invoke19_go_in = ~(pd51_out | invoke19_done_out) & par0_go_out;
    assign invoke1_done_in = me2_done;
    assign invoke1_go_in = ~(pd33_out | invoke1_done_out) & par0_go_out;
    assign invoke20_done_in = me21_done;
    assign invoke20_go_in = ~(pd52_out | invoke20_done_out) & par0_go_out;
    assign invoke21_done_in = me22_done;
    assign invoke21_go_in = ~(pd53_out | invoke21_done_out) & par0_go_out;
    assign invoke22_done_in = me23_done;
    assign invoke22_go_in = ~(pd54_out | invoke22_done_out) & par0_go_out;
    assign invoke23_done_in = me24_done;
    assign invoke23_go_in = ~(pd55_out | invoke23_done_out) & par0_go_out;
    assign invoke24_done_in = me25_done;
    assign invoke24_go_in = ~(pd56_out | invoke24_done_out) & par0_go_out;
    assign invoke25_done_in = me26_done;
    assign invoke25_go_in = ~(pd57_out | invoke25_done_out) & par0_go_out;
    assign invoke26_done_in = me27_done;
    assign invoke26_go_in = ~(pd58_out | invoke26_done_out) & par0_go_out;
    assign invoke27_done_in = me28_done;
    assign invoke27_go_in = ~(pd59_out | invoke27_done_out) & par0_go_out;
    assign invoke28_done_in = me29_done;
    assign invoke28_go_in = ~(pd60_out | invoke28_done_out) & par0_go_out;
    assign invoke29_done_in = me30_done;
    assign invoke29_go_in = ~(pd61_out | invoke29_done_out) & par0_go_out;
    assign invoke2_done_in = me3_done;
    assign invoke2_go_in = ~(pd34_out | invoke2_done_out) & par0_go_out;
    assign invoke30_done_in = me31_done;
    assign invoke30_go_in = ~(pd62_out | invoke30_done_out) & par0_go_out;
    assign invoke31_done_in = ce00_done;
    assign invoke31_go_in = ~(pd63_out | invoke31_done_out) & par1_go_out;
    assign invoke32_done_in = ce01_done;
    assign invoke32_go_in = ~(pd64_out | invoke32_done_out) & par1_go_out;
    assign invoke33_done_in = ce02_done;
    assign invoke33_go_in = ~(pd65_out | invoke33_done_out) & par1_go_out;
    assign invoke34_done_in = ce03_done;
    assign invoke34_go_in = ~(pd66_out | invoke34_done_out) & par1_go_out;
    assign invoke35_done_in = ce04_done;
    assign invoke35_go_in = ~(pd67_out | invoke35_done_out) & par1_go_out;
    assign invoke36_done_in = ce05_done;
    assign invoke36_go_in = ~(pd68_out | invoke36_done_out) & par1_go_out;
    assign invoke37_done_in = ce06_done;
    assign invoke37_go_in = ~(pd69_out | invoke37_done_out) & par1_go_out;
    assign invoke38_done_in = ce07_done;
    assign invoke38_go_in = ~(pd70_out | invoke38_done_out) & par1_go_out;
    assign invoke39_done_in = ce08_done;
    assign invoke39_go_in = ~(pd71_out | invoke39_done_out) & par1_go_out;
    assign invoke3_done_in = me4_done;
    assign invoke3_go_in = ~(pd35_out | invoke3_done_out) & par0_go_out;
    assign invoke40_done_in = ce09_done;
    assign invoke40_go_in = ~(pd72_out | invoke40_done_out) & par1_go_out;
    assign invoke41_done_in = ce010_done;
    assign invoke41_go_in = ~(pd73_out | invoke41_done_out) & par1_go_out;
    assign invoke42_done_in = ce011_done;
    assign invoke42_go_in = ~(pd74_out | invoke42_done_out) & par1_go_out;
    assign invoke43_done_in = ce012_done;
    assign invoke43_go_in = ~(pd75_out | invoke43_done_out) & par1_go_out;
    assign invoke44_done_in = ce013_done;
    assign invoke44_go_in = ~(pd76_out | invoke44_done_out) & par1_go_out;
    assign invoke45_done_in = ce014_done;
    assign invoke45_go_in = ~(pd77_out | invoke45_done_out) & par1_go_out;
    assign invoke46_done_in = ce015_done;
    assign invoke46_go_in = ~(pd78_out | invoke46_done_out) & par1_go_out;
    assign invoke47_done_in = ce10_done;
    assign invoke47_go_in = ~(pd79_out | invoke47_done_out) & par2_go_out;
    assign invoke48_done_in = ce11_done;
    assign invoke48_go_in = ~(pd80_out | invoke48_done_out) & par2_go_out;
    assign invoke49_done_in = ce12_done;
    assign invoke49_go_in = ~(pd81_out | invoke49_done_out) & par2_go_out;
    assign invoke4_done_in = me5_done;
    assign invoke4_go_in = ~(pd36_out | invoke4_done_out) & par0_go_out;
    assign invoke50_done_in = ce13_done;
    assign invoke50_go_in = ~(pd82_out | invoke50_done_out) & par2_go_out;
    assign invoke51_done_in = ce14_done;
    assign invoke51_go_in = ~(pd83_out | invoke51_done_out) & par2_go_out;
    assign invoke52_done_in = ce15_done;
    assign invoke52_go_in = ~(pd84_out | invoke52_done_out) & par2_go_out;
    assign invoke53_done_in = ce16_done;
    assign invoke53_go_in = ~(pd85_out | invoke53_done_out) & par2_go_out;
    assign invoke54_done_in = ce17_done;
    assign invoke54_go_in = ~(pd86_out | invoke54_done_out) & par2_go_out;
    assign invoke55_done_in = ce20_done;
    assign invoke55_go_in = ~(pd87_out | invoke55_done_out) & par3_go_out;
    assign invoke56_done_in = ce21_done;
    assign invoke56_go_in = ~(pd88_out | invoke56_done_out) & par3_go_out;
    assign invoke57_done_in = ce22_done;
    assign invoke57_go_in = ~(pd89_out | invoke57_done_out) & par3_go_out;
    assign invoke58_done_in = ce23_done;
    assign invoke58_go_in = ~(pd90_out | invoke58_done_out) & par3_go_out;
    assign invoke59_done_in = ce30_done;
    assign invoke59_go_in = ~(pd91_out | invoke59_done_out) & par4_go_out;
    assign invoke5_done_in = me6_done;
    assign invoke5_go_in = ~(pd37_out | invoke5_done_out) & par0_go_out;
    assign invoke60_done_in = ce31_done;
    assign invoke60_go_in = ~(pd92_out | invoke60_done_out) & par4_go_out;
    assign invoke61_done_in = ce40_done;
    assign invoke61_go_in = ~invoke61_done_out & fsm32_out == 4'd6 & tdcc32_go_out;
    assign invoke6_done_in = me7_done;
    assign invoke6_go_in = ~(pd38_out | invoke6_done_out) & par0_go_out;
    assign invoke7_done_in = me8_done;
    assign invoke7_go_in = ~(pd39_out | invoke7_done_out) & par0_go_out;
    assign invoke8_done_in = me9_done;
    assign invoke8_go_in = ~(pd40_out | invoke8_done_out) & par0_go_out;
    assign invoke9_done_in = me10_done;
    assign invoke9_go_in = ~(pd41_out | invoke9_done_out) & par0_go_out;
    assign invoke_done_in = me0_done;
    assign invoke_go_in = ~(pd31_out | invoke_done_out) & par0_go_out;
    assign is_index0_left =
     find_write_index_go_out ? 5'd0 : 5'd0;
    assign is_index0_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index1_left =
     find_write_index_go_out ? 5'd1 : 5'd0;
    assign is_index1_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index10_left =
     find_write_index_go_out ? 5'd10 : 5'd0;
    assign is_index10_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index11_left =
     find_write_index_go_out ? 5'd11 : 5'd0;
    assign is_index11_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index12_left =
     find_write_index_go_out ? 5'd12 : 5'd0;
    assign is_index12_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index13_left =
     find_write_index_go_out ? 5'd13 : 5'd0;
    assign is_index13_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index14_left =
     find_write_index_go_out ? 5'd14 : 5'd0;
    assign is_index14_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index15_left =
     find_write_index_go_out ? 5'd15 : 5'd0;
    assign is_index15_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index16_left =
     find_write_index_go_out ? 5'd16 : 5'd0;
    assign is_index16_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index17_left =
     find_write_index_go_out ? 5'd17 : 5'd0;
    assign is_index17_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index18_left =
     find_write_index_go_out ? 5'd18 : 5'd0;
    assign is_index18_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index19_left =
     find_write_index_go_out ? 5'd19 : 5'd0;
    assign is_index19_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index2_left =
     find_write_index_go_out ? 5'd2 : 5'd0;
    assign is_index2_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index20_left =
     find_write_index_go_out ? 5'd20 : 5'd0;
    assign is_index20_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index21_left =
     find_write_index_go_out ? 5'd21 : 5'd0;
    assign is_index21_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index22_left =
     find_write_index_go_out ? 5'd22 : 5'd0;
    assign is_index22_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index23_left =
     find_write_index_go_out ? 5'd23 : 5'd0;
    assign is_index23_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index24_left =
     find_write_index_go_out ? 5'd24 : 5'd0;
    assign is_index24_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index25_left =
     find_write_index_go_out ? 5'd25 : 5'd0;
    assign is_index25_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index26_left =
     find_write_index_go_out ? 5'd26 : 5'd0;
    assign is_index26_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index27_left =
     find_write_index_go_out ? 5'd27 : 5'd0;
    assign is_index27_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index28_left =
     find_write_index_go_out ? 5'd28 : 5'd0;
    assign is_index28_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index29_left =
     find_write_index_go_out ? 5'd29 : 5'd0;
    assign is_index29_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index3_left =
     find_write_index_go_out ? 5'd3 : 5'd0;
    assign is_index3_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index30_left =
     find_write_index_go_out ? 5'd30 : 5'd0;
    assign is_index30_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index31_left =
     find_write_index_go_out ? 5'd31 : 5'd0;
    assign is_index31_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index4_left =
     find_write_index_go_out ? 5'd4 : 5'd0;
    assign is_index4_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index5_left =
     find_write_index_go_out ? 5'd5 : 5'd0;
    assign is_index5_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index6_left =
     find_write_index_go_out ? 5'd6 : 5'd0;
    assign is_index6_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index7_left =
     find_write_index_go_out ? 5'd7 : 5'd0;
    assign is_index7_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index8_left =
     find_write_index_go_out ? 5'd8 : 5'd0;
    assign is_index8_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_index9_left =
     find_write_index_go_out ? 5'd9 : 5'd0;
    assign is_index9_right =
     find_write_index_go_out ? write_index : 5'd0;
    assign is_length_zero0_done_in = comb_reg1_done;
    assign is_length_zero0_go_in = ~is_length_zero0_done_out & fsm31_out == 3'd1 & tdcc31_go_out;
    assign l0_clk = clk;
    assign l0_in =
     write0_go_out ? slice_out : 5'd0;
    assign l0_reset = reset;
    assign l0_write_en =
     write0_go_out ? write_en : 1'd0;
    assign l1_clk = clk;
    assign l1_in =
     write1_go_out ? slice_out : 5'd0;
    assign l1_reset = reset;
    assign l1_write_en =
     write1_go_out ? write_en : 1'd0;
    assign l10_clk = clk;
    assign l10_in =
     write10_go_out ? slice_out : 5'd0;
    assign l10_reset = reset;
    assign l10_write_en =
     write10_go_out ? write_en : 1'd0;
    assign l11_clk = clk;
    assign l11_in =
     write11_go_out ? slice_out : 5'd0;
    assign l11_reset = reset;
    assign l11_write_en =
     write11_go_out ? write_en : 1'd0;
    assign l12_clk = clk;
    assign l12_in =
     write12_go_out ? slice_out : 5'd0;
    assign l12_reset = reset;
    assign l12_write_en =
     write12_go_out ? write_en : 1'd0;
    assign l13_clk = clk;
    assign l13_in =
     write13_go_out ? slice_out : 5'd0;
    assign l13_reset = reset;
    assign l13_write_en =
     write13_go_out ? write_en : 1'd0;
    assign l14_clk = clk;
    assign l14_in =
     write14_go_out ? slice_out : 5'd0;
    assign l14_reset = reset;
    assign l14_write_en =
     write14_go_out ? write_en : 1'd0;
    assign l15_clk = clk;
    assign l15_in =
     write15_go_out ? slice_out : 5'd0;
    assign l15_reset = reset;
    assign l15_write_en =
     write15_go_out ? write_en : 1'd0;
    assign l16_clk = clk;
    assign l16_in =
     write16_go_out ? slice_out : 5'd0;
    assign l16_reset = reset;
    assign l16_write_en =
     write16_go_out ? write_en : 1'd0;
    assign l17_clk = clk;
    assign l17_in =
     write17_go_out ? slice_out : 5'd0;
    assign l17_reset = reset;
    assign l17_write_en =
     write17_go_out ? write_en : 1'd0;
    assign l18_clk = clk;
    assign l18_in =
     write18_go_out ? slice_out : 5'd0;
    assign l18_reset = reset;
    assign l18_write_en =
     write18_go_out ? write_en : 1'd0;
    assign l19_clk = clk;
    assign l19_in =
     write19_go_out ? slice_out : 5'd0;
    assign l19_reset = reset;
    assign l19_write_en =
     write19_go_out ? write_en : 1'd0;
    assign l2_clk = clk;
    assign l2_in =
     write2_go_out ? slice_out : 5'd0;
    assign l2_reset = reset;
    assign l2_write_en =
     write2_go_out ? write_en : 1'd0;
    assign l20_clk = clk;
    assign l20_in =
     write20_go_out ? slice_out : 5'd0;
    assign l20_reset = reset;
    assign l20_write_en =
     write20_go_out ? write_en : 1'd0;
    assign l21_clk = clk;
    assign l21_in =
     write21_go_out ? slice_out : 5'd0;
    assign l21_reset = reset;
    assign l21_write_en =
     write21_go_out ? write_en : 1'd0;
    assign l22_clk = clk;
    assign l22_in =
     write22_go_out ? slice_out : 5'd0;
    assign l22_reset = reset;
    assign l22_write_en =
     write22_go_out ? write_en : 1'd0;
    assign l23_clk = clk;
    assign l23_in =
     write23_go_out ? slice_out : 5'd0;
    assign l23_reset = reset;
    assign l23_write_en =
     write23_go_out ? write_en : 1'd0;
    assign l24_clk = clk;
    assign l24_in =
     write24_go_out ? slice_out : 5'd0;
    assign l24_reset = reset;
    assign l24_write_en =
     write24_go_out ? write_en : 1'd0;
    assign l25_clk = clk;
    assign l25_in =
     write25_go_out ? slice_out : 5'd0;
    assign l25_reset = reset;
    assign l25_write_en =
     write25_go_out ? write_en : 1'd0;
    assign l26_clk = clk;
    assign l26_in =
     write26_go_out ? slice_out : 5'd0;
    assign l26_reset = reset;
    assign l26_write_en =
     write26_go_out ? write_en : 1'd0;
    assign l27_clk = clk;
    assign l27_in =
     write27_go_out ? slice_out : 5'd0;
    assign l27_reset = reset;
    assign l27_write_en =
     write27_go_out ? write_en : 1'd0;
    assign l28_clk = clk;
    assign l28_in =
     write28_go_out ? slice_out : 5'd0;
    assign l28_reset = reset;
    assign l28_write_en =
     write28_go_out ? write_en : 1'd0;
    assign l29_clk = clk;
    assign l29_in =
     write29_go_out ? slice_out : 5'd0;
    assign l29_reset = reset;
    assign l29_write_en =
     write29_go_out ? write_en : 1'd0;
    assign l3_clk = clk;
    assign l3_in =
     write3_go_out ? slice_out : 5'd0;
    assign l3_reset = reset;
    assign l3_write_en =
     write3_go_out ? write_en : 1'd0;
    assign l30_clk = clk;
    assign l30_in =
     write30_go_out ? slice_out : 5'd0;
    assign l30_reset = reset;
    assign l30_write_en =
     write30_go_out ? write_en : 1'd0;
    assign l31_clk = clk;
    assign l31_in =
     write31_go_out ? slice_out : 5'd0;
    assign l31_reset = reset;
    assign l31_write_en =
     write31_go_out ? write_en : 1'd0;
    assign l4_clk = clk;
    assign l4_in =
     write4_go_out ? slice_out : 5'd0;
    assign l4_reset = reset;
    assign l4_write_en =
     write4_go_out ? write_en : 1'd0;
    assign l5_clk = clk;
    assign l5_in =
     write5_go_out ? slice_out : 5'd0;
    assign l5_reset = reset;
    assign l5_write_en =
     write5_go_out ? write_en : 1'd0;
    assign l6_clk = clk;
    assign l6_in =
     write6_go_out ? slice_out : 5'd0;
    assign l6_reset = reset;
    assign l6_write_en =
     write6_go_out ? write_en : 1'd0;
    assign l7_clk = clk;
    assign l7_in =
     write7_go_out ? slice_out : 5'd0;
    assign l7_reset = reset;
    assign l7_write_en =
     write7_go_out ? write_en : 1'd0;
    assign l8_clk = clk;
    assign l8_in =
     write8_go_out ? slice_out : 5'd0;
    assign l8_reset = reset;
    assign l8_write_en =
     write8_go_out ? write_en : 1'd0;
    assign l9_clk = clk;
    assign l9_in =
     write9_go_out ? slice_out : 5'd0;
    assign l9_reset = reset;
    assign l9_write_en =
     write9_go_out ? write_en : 1'd0;
    assign me0_clk = clk;
    assign me0_go = invoke_go_out;
    assign me0_in =
     invoke_go_out ? in : 32'd0;
    assign me0_length =
     invoke_go_out ? l0_out : 5'd0;
    assign me0_prefix =
     invoke_go_out ? p0_out : 32'd0;
    assign me0_reset = reset;
    assign me1_clk = clk;
    assign me1_go = invoke0_go_out;
    assign me1_in =
     invoke0_go_out ? in : 32'd0;
    assign me1_length =
     invoke0_go_out ? l1_out : 5'd0;
    assign me1_prefix =
     invoke0_go_out ? p1_out : 32'd0;
    assign me1_reset = reset;
    assign me10_clk = clk;
    assign me10_go = invoke9_go_out;
    assign me10_in =
     invoke9_go_out ? in : 32'd0;
    assign me10_length =
     invoke9_go_out ? l10_out : 5'd0;
    assign me10_prefix =
     invoke9_go_out ? p10_out : 32'd0;
    assign me10_reset = reset;
    assign me11_clk = clk;
    assign me11_go = invoke10_go_out;
    assign me11_in =
     invoke10_go_out ? in : 32'd0;
    assign me11_length =
     invoke10_go_out ? l11_out : 5'd0;
    assign me11_prefix =
     invoke10_go_out ? p11_out : 32'd0;
    assign me11_reset = reset;
    assign me12_clk = clk;
    assign me12_go = invoke11_go_out;
    assign me12_in =
     invoke11_go_out ? in : 32'd0;
    assign me12_length =
     invoke11_go_out ? l12_out : 5'd0;
    assign me12_prefix =
     invoke11_go_out ? p12_out : 32'd0;
    assign me12_reset = reset;
    assign me13_clk = clk;
    assign me13_go = invoke12_go_out;
    assign me13_in =
     invoke12_go_out ? in : 32'd0;
    assign me13_length =
     invoke12_go_out ? l13_out : 5'd0;
    assign me13_prefix =
     invoke12_go_out ? p13_out : 32'd0;
    assign me13_reset = reset;
    assign me14_clk = clk;
    assign me14_go = invoke13_go_out;
    assign me14_in =
     invoke13_go_out ? in : 32'd0;
    assign me14_length =
     invoke13_go_out ? l14_out : 5'd0;
    assign me14_prefix =
     invoke13_go_out ? p14_out : 32'd0;
    assign me14_reset = reset;
    assign me15_clk = clk;
    assign me15_go = invoke14_go_out;
    assign me15_in =
     invoke14_go_out ? in : 32'd0;
    assign me15_length =
     invoke14_go_out ? l15_out : 5'd0;
    assign me15_prefix =
     invoke14_go_out ? p15_out : 32'd0;
    assign me15_reset = reset;
    assign me16_clk = clk;
    assign me16_go = invoke15_go_out;
    assign me16_in =
     invoke15_go_out ? in : 32'd0;
    assign me16_length =
     invoke15_go_out ? l16_out : 5'd0;
    assign me16_prefix =
     invoke15_go_out ? p16_out : 32'd0;
    assign me16_reset = reset;
    assign me17_clk = clk;
    assign me17_go = invoke16_go_out;
    assign me17_in =
     invoke16_go_out ? in : 32'd0;
    assign me17_length =
     invoke16_go_out ? l17_out : 5'd0;
    assign me17_prefix =
     invoke16_go_out ? p17_out : 32'd0;
    assign me17_reset = reset;
    assign me18_clk = clk;
    assign me18_go = invoke17_go_out;
    assign me18_in =
     invoke17_go_out ? in : 32'd0;
    assign me18_length =
     invoke17_go_out ? l18_out : 5'd0;
    assign me18_prefix =
     invoke17_go_out ? p18_out : 32'd0;
    assign me18_reset = reset;
    assign me19_clk = clk;
    assign me19_go = invoke18_go_out;
    assign me19_in =
     invoke18_go_out ? in : 32'd0;
    assign me19_length =
     invoke18_go_out ? l19_out : 5'd0;
    assign me19_prefix =
     invoke18_go_out ? p19_out : 32'd0;
    assign me19_reset = reset;
    assign me2_clk = clk;
    assign me2_go = invoke1_go_out;
    assign me2_in =
     invoke1_go_out ? in : 32'd0;
    assign me2_length =
     invoke1_go_out ? l2_out : 5'd0;
    assign me2_prefix =
     invoke1_go_out ? p2_out : 32'd0;
    assign me2_reset = reset;
    assign me20_clk = clk;
    assign me20_go = invoke19_go_out;
    assign me20_in =
     invoke19_go_out ? in : 32'd0;
    assign me20_length =
     invoke19_go_out ? l20_out : 5'd0;
    assign me20_prefix =
     invoke19_go_out ? p20_out : 32'd0;
    assign me20_reset = reset;
    assign me21_clk = clk;
    assign me21_go = invoke20_go_out;
    assign me21_in =
     invoke20_go_out ? in : 32'd0;
    assign me21_length =
     invoke20_go_out ? l21_out : 5'd0;
    assign me21_prefix =
     invoke20_go_out ? p21_out : 32'd0;
    assign me21_reset = reset;
    assign me22_clk = clk;
    assign me22_go = invoke21_go_out;
    assign me22_in =
     invoke21_go_out ? in : 32'd0;
    assign me22_length =
     invoke21_go_out ? l22_out : 5'd0;
    assign me22_prefix =
     invoke21_go_out ? p22_out : 32'd0;
    assign me22_reset = reset;
    assign me23_clk = clk;
    assign me23_go = invoke22_go_out;
    assign me23_in =
     invoke22_go_out ? in : 32'd0;
    assign me23_length =
     invoke22_go_out ? l23_out : 5'd0;
    assign me23_prefix =
     invoke22_go_out ? p23_out : 32'd0;
    assign me23_reset = reset;
    assign me24_clk = clk;
    assign me24_go = invoke23_go_out;
    assign me24_in =
     invoke23_go_out ? in : 32'd0;
    assign me24_length =
     invoke23_go_out ? l24_out : 5'd0;
    assign me24_prefix =
     invoke23_go_out ? p24_out : 32'd0;
    assign me24_reset = reset;
    assign me25_clk = clk;
    assign me25_go = invoke24_go_out;
    assign me25_in =
     invoke24_go_out ? in : 32'd0;
    assign me25_length =
     invoke24_go_out ? l25_out : 5'd0;
    assign me25_prefix =
     invoke24_go_out ? p25_out : 32'd0;
    assign me25_reset = reset;
    assign me26_clk = clk;
    assign me26_go = invoke25_go_out;
    assign me26_in =
     invoke25_go_out ? in : 32'd0;
    assign me26_length =
     invoke25_go_out ? l26_out : 5'd0;
    assign me26_prefix =
     invoke25_go_out ? p26_out : 32'd0;
    assign me26_reset = reset;
    assign me27_clk = clk;
    assign me27_go = invoke26_go_out;
    assign me27_in =
     invoke26_go_out ? in : 32'd0;
    assign me27_length =
     invoke26_go_out ? l27_out : 5'd0;
    assign me27_prefix =
     invoke26_go_out ? p27_out : 32'd0;
    assign me27_reset = reset;
    assign me28_clk = clk;
    assign me28_go = invoke27_go_out;
    assign me28_in =
     invoke27_go_out ? in : 32'd0;
    assign me28_length =
     invoke27_go_out ? l28_out : 5'd0;
    assign me28_prefix =
     invoke27_go_out ? p28_out : 32'd0;
    assign me28_reset = reset;
    assign me29_clk = clk;
    assign me29_go = invoke28_go_out;
    assign me29_in =
     invoke28_go_out ? in : 32'd0;
    assign me29_length =
     invoke28_go_out ? l29_out : 5'd0;
    assign me29_prefix =
     invoke28_go_out ? p29_out : 32'd0;
    assign me29_reset = reset;
    assign me3_clk = clk;
    assign me3_go = invoke2_go_out;
    assign me3_in =
     invoke2_go_out ? in : 32'd0;
    assign me3_length =
     invoke2_go_out ? l3_out : 5'd0;
    assign me3_prefix =
     invoke2_go_out ? p3_out : 32'd0;
    assign me3_reset = reset;
    assign me30_clk = clk;
    assign me30_go = invoke29_go_out;
    assign me30_in =
     invoke29_go_out ? in : 32'd0;
    assign me30_length =
     invoke29_go_out ? l30_out : 5'd0;
    assign me30_prefix =
     invoke29_go_out ? p30_out : 32'd0;
    assign me30_reset = reset;
    assign me31_clk = clk;
    assign me31_go = invoke30_go_out;
    assign me31_in =
     invoke30_go_out ? in : 32'd0;
    assign me31_length =
     invoke30_go_out ? l31_out : 5'd0;
    assign me31_prefix =
     invoke30_go_out ? p31_out : 32'd0;
    assign me31_reset = reset;
    assign me4_clk = clk;
    assign me4_go = invoke3_go_out;
    assign me4_in =
     invoke3_go_out ? in : 32'd0;
    assign me4_length =
     invoke3_go_out ? l4_out : 5'd0;
    assign me4_prefix =
     invoke3_go_out ? p4_out : 32'd0;
    assign me4_reset = reset;
    assign me5_clk = clk;
    assign me5_go = invoke4_go_out;
    assign me5_in =
     invoke4_go_out ? in : 32'd0;
    assign me5_length =
     invoke4_go_out ? l5_out : 5'd0;
    assign me5_prefix =
     invoke4_go_out ? p5_out : 32'd0;
    assign me5_reset = reset;
    assign me6_clk = clk;
    assign me6_go = invoke5_go_out;
    assign me6_in =
     invoke5_go_out ? in : 32'd0;
    assign me6_length =
     invoke5_go_out ? l6_out : 5'd0;
    assign me6_prefix =
     invoke5_go_out ? p6_out : 32'd0;
    assign me6_reset = reset;
    assign me7_clk = clk;
    assign me7_go = invoke6_go_out;
    assign me7_in =
     invoke6_go_out ? in : 32'd0;
    assign me7_length =
     invoke6_go_out ? l7_out : 5'd0;
    assign me7_prefix =
     invoke6_go_out ? p7_out : 32'd0;
    assign me7_reset = reset;
    assign me8_clk = clk;
    assign me8_go = invoke7_go_out;
    assign me8_in =
     invoke7_go_out ? in : 32'd0;
    assign me8_length =
     invoke7_go_out ? l8_out : 5'd0;
    assign me8_prefix =
     invoke7_go_out ? p8_out : 32'd0;
    assign me8_reset = reset;
    assign me9_clk = clk;
    assign me9_go = invoke8_go_out;
    assign me9_in =
     invoke8_go_out ? in : 32'd0;
    assign me9_length =
     invoke8_go_out ? l9_out : 5'd0;
    assign me9_prefix =
     invoke8_go_out ? p9_out : 32'd0;
    assign me9_reset = reset;
    assign out_clk = clk;
    assign out_in =
     save_index_go_out ? ce40_addrX :
     default_to_zero_length_index_go_out ? zero_index_out : 5'd0;
    assign out_reset = reset;
    assign out_write_en = default_to_zero_length_index_go_out | save_index_go_out;
    assign p0_clk = clk;
    assign p0_in =
     write0_go_out ? in : 32'd0;
    assign p0_reset = reset;
    assign p0_write_en =
     write0_go_out ? write_en : 1'd0;
    assign p1_clk = clk;
    assign p1_in =
     write1_go_out ? in : 32'd0;
    assign p1_reset = reset;
    assign p1_write_en =
     write1_go_out ? write_en : 1'd0;
    assign p10_clk = clk;
    assign p10_in =
     write10_go_out ? in : 32'd0;
    assign p10_reset = reset;
    assign p10_write_en =
     write10_go_out ? write_en : 1'd0;
    assign p11_clk = clk;
    assign p11_in =
     write11_go_out ? in : 32'd0;
    assign p11_reset = reset;
    assign p11_write_en =
     write11_go_out ? write_en : 1'd0;
    assign p12_clk = clk;
    assign p12_in =
     write12_go_out ? in : 32'd0;
    assign p12_reset = reset;
    assign p12_write_en =
     write12_go_out ? write_en : 1'd0;
    assign p13_clk = clk;
    assign p13_in =
     write13_go_out ? in : 32'd0;
    assign p13_reset = reset;
    assign p13_write_en =
     write13_go_out ? write_en : 1'd0;
    assign p14_clk = clk;
    assign p14_in =
     write14_go_out ? in : 32'd0;
    assign p14_reset = reset;
    assign p14_write_en =
     write14_go_out ? write_en : 1'd0;
    assign p15_clk = clk;
    assign p15_in =
     write15_go_out ? in : 32'd0;
    assign p15_reset = reset;
    assign p15_write_en =
     write15_go_out ? write_en : 1'd0;
    assign p16_clk = clk;
    assign p16_in =
     write16_go_out ? in : 32'd0;
    assign p16_reset = reset;
    assign p16_write_en =
     write16_go_out ? write_en : 1'd0;
    assign p17_clk = clk;
    assign p17_in =
     write17_go_out ? in : 32'd0;
    assign p17_reset = reset;
    assign p17_write_en =
     write17_go_out ? write_en : 1'd0;
    assign p18_clk = clk;
    assign p18_in =
     write18_go_out ? in : 32'd0;
    assign p18_reset = reset;
    assign p18_write_en =
     write18_go_out ? write_en : 1'd0;
    assign p19_clk = clk;
    assign p19_in =
     write19_go_out ? in : 32'd0;
    assign p19_reset = reset;
    assign p19_write_en =
     write19_go_out ? write_en : 1'd0;
    assign p2_clk = clk;
    assign p2_in =
     write2_go_out ? in : 32'd0;
    assign p2_reset = reset;
    assign p2_write_en =
     write2_go_out ? write_en : 1'd0;
    assign p20_clk = clk;
    assign p20_in =
     write20_go_out ? in : 32'd0;
    assign p20_reset = reset;
    assign p20_write_en =
     write20_go_out ? write_en : 1'd0;
    assign p21_clk = clk;
    assign p21_in =
     write21_go_out ? in : 32'd0;
    assign p21_reset = reset;
    assign p21_write_en =
     write21_go_out ? write_en : 1'd0;
    assign p22_clk = clk;
    assign p22_in =
     write22_go_out ? in : 32'd0;
    assign p22_reset = reset;
    assign p22_write_en =
     write22_go_out ? write_en : 1'd0;
    assign p23_clk = clk;
    assign p23_in =
     write23_go_out ? in : 32'd0;
    assign p23_reset = reset;
    assign p23_write_en =
     write23_go_out ? write_en : 1'd0;
    assign p24_clk = clk;
    assign p24_in =
     write24_go_out ? in : 32'd0;
    assign p24_reset = reset;
    assign p24_write_en =
     write24_go_out ? write_en : 1'd0;
    assign p25_clk = clk;
    assign p25_in =
     write25_go_out ? in : 32'd0;
    assign p25_reset = reset;
    assign p25_write_en =
     write25_go_out ? write_en : 1'd0;
    assign p26_clk = clk;
    assign p26_in =
     write26_go_out ? in : 32'd0;
    assign p26_reset = reset;
    assign p26_write_en =
     write26_go_out ? write_en : 1'd0;
    assign p27_clk = clk;
    assign p27_in =
     write27_go_out ? in : 32'd0;
    assign p27_reset = reset;
    assign p27_write_en =
     write27_go_out ? write_en : 1'd0;
    assign p28_clk = clk;
    assign p28_in =
     write28_go_out ? in : 32'd0;
    assign p28_reset = reset;
    assign p28_write_en =
     write28_go_out ? write_en : 1'd0;
    assign p29_clk = clk;
    assign p29_in =
     write29_go_out ? in : 32'd0;
    assign p29_reset = reset;
    assign p29_write_en =
     write29_go_out ? write_en : 1'd0;
    assign p3_clk = clk;
    assign p3_in =
     write3_go_out ? in : 32'd0;
    assign p3_reset = reset;
    assign p3_write_en =
     write3_go_out ? write_en : 1'd0;
    assign p30_clk = clk;
    assign p30_in =
     write30_go_out ? in : 32'd0;
    assign p30_reset = reset;
    assign p30_write_en =
     write30_go_out ? write_en : 1'd0;
    assign p31_clk = clk;
    assign p31_in =
     write31_go_out ? in : 32'd0;
    assign p31_reset = reset;
    assign p31_write_en =
     write31_go_out ? write_en : 1'd0;
    assign p4_clk = clk;
    assign p4_in =
     write4_go_out ? in : 32'd0;
    assign p4_reset = reset;
    assign p4_write_en =
     write4_go_out ? write_en : 1'd0;
    assign p5_clk = clk;
    assign p5_in =
     write5_go_out ? in : 32'd0;
    assign p5_reset = reset;
    assign p5_write_en =
     write5_go_out ? write_en : 1'd0;
    assign p6_clk = clk;
    assign p6_in =
     write6_go_out ? in : 32'd0;
    assign p6_reset = reset;
    assign p6_write_en =
     write6_go_out ? write_en : 1'd0;
    assign p7_clk = clk;
    assign p7_in =
     write7_go_out ? in : 32'd0;
    assign p7_reset = reset;
    assign p7_write_en =
     write7_go_out ? write_en : 1'd0;
    assign p8_clk = clk;
    assign p8_in =
     write8_go_out ? in : 32'd0;
    assign p8_reset = reset;
    assign p8_write_en =
     write8_go_out ? write_en : 1'd0;
    assign p9_clk = clk;
    assign p9_in =
     write9_go_out ? in : 32'd0;
    assign p9_reset = reset;
    assign p9_write_en =
     write9_go_out ? write_en : 1'd0;
    assign par0_done_in = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out;
    assign par0_go_in = ~par0_done_out & fsm32_out == 4'd1 & tdcc32_go_out;
    assign par1_done_in = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out;
    assign par1_go_in = ~par1_done_out & fsm32_out == 4'd2 & tdcc32_go_out;
    assign par2_done_in = pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out;
    assign par2_go_in = ~par2_done_out & fsm32_out == 4'd3 & tdcc32_go_out;
    assign par3_done_in = pd87_out & pd88_out & pd89_out & pd90_out;
    assign par3_go_in = ~par3_done_out & fsm32_out == 4'd4 & tdcc32_go_out;
    assign par4_done_in = pd91_out & pd92_out;
    assign par4_go_in = ~par4_done_out & fsm32_out == 4'd5 & tdcc32_go_out;
    assign par5_done_in = pd93_out & pd94_out;
    assign par5_go_in = ~par5_done_out & fsm33_out == 1'd0 & tdcc33_go_out;
    assign par_done_in = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out;
    assign par_go_in = ~par_done_out & fsm31_out == 3'd4 & tdcc31_go_out;
    assign pd_clk = clk;
    assign pd_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd_reset = reset;
    assign pd_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc_done_out & par_go_out;
    assign pd0_clk = clk;
    assign pd0_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc0_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd0_reset = reset;
    assign pd0_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc0_done_out & par_go_out;
    assign pd1_clk = clk;
    assign pd1_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc1_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd1_reset = reset;
    assign pd1_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc1_done_out & par_go_out;
    assign pd10_clk = clk;
    assign pd10_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc10_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd10_reset = reset;
    assign pd10_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc10_done_out & par_go_out;
    assign pd11_clk = clk;
    assign pd11_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc11_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd11_reset = reset;
    assign pd11_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc11_done_out & par_go_out;
    assign pd12_clk = clk;
    assign pd12_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc12_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd12_reset = reset;
    assign pd12_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc12_done_out & par_go_out;
    assign pd13_clk = clk;
    assign pd13_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc13_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd13_reset = reset;
    assign pd13_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc13_done_out & par_go_out;
    assign pd14_clk = clk;
    assign pd14_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc14_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd14_reset = reset;
    assign pd14_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc14_done_out & par_go_out;
    assign pd15_clk = clk;
    assign pd15_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc15_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd15_reset = reset;
    assign pd15_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc15_done_out & par_go_out;
    assign pd16_clk = clk;
    assign pd16_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc16_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd16_reset = reset;
    assign pd16_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc16_done_out & par_go_out;
    assign pd17_clk = clk;
    assign pd17_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc17_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd17_reset = reset;
    assign pd17_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc17_done_out & par_go_out;
    assign pd18_clk = clk;
    assign pd18_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc18_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd18_reset = reset;
    assign pd18_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc18_done_out & par_go_out;
    assign pd19_clk = clk;
    assign pd19_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc19_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd19_reset = reset;
    assign pd19_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc19_done_out & par_go_out;
    assign pd2_clk = clk;
    assign pd2_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc2_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd2_reset = reset;
    assign pd2_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc2_done_out & par_go_out;
    assign pd20_clk = clk;
    assign pd20_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc20_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd20_reset = reset;
    assign pd20_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc20_done_out & par_go_out;
    assign pd21_clk = clk;
    assign pd21_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc21_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd21_reset = reset;
    assign pd21_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc21_done_out & par_go_out;
    assign pd22_clk = clk;
    assign pd22_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc22_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd22_reset = reset;
    assign pd22_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc22_done_out & par_go_out;
    assign pd23_clk = clk;
    assign pd23_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc23_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd23_reset = reset;
    assign pd23_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc23_done_out & par_go_out;
    assign pd24_clk = clk;
    assign pd24_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc24_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd24_reset = reset;
    assign pd24_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc24_done_out & par_go_out;
    assign pd25_clk = clk;
    assign pd25_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc25_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd25_reset = reset;
    assign pd25_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc25_done_out & par_go_out;
    assign pd26_clk = clk;
    assign pd26_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc26_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd26_reset = reset;
    assign pd26_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc26_done_out & par_go_out;
    assign pd27_clk = clk;
    assign pd27_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc27_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd27_reset = reset;
    assign pd27_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc27_done_out & par_go_out;
    assign pd28_clk = clk;
    assign pd28_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc28_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd28_reset = reset;
    assign pd28_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc28_done_out & par_go_out;
    assign pd29_clk = clk;
    assign pd29_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc29_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd29_reset = reset;
    assign pd29_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc29_done_out & par_go_out;
    assign pd3_clk = clk;
    assign pd3_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc3_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd3_reset = reset;
    assign pd3_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc3_done_out & par_go_out;
    assign pd30_clk = clk;
    assign pd30_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc30_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd30_reset = reset;
    assign pd30_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc30_done_out & par_go_out;
    assign pd31_clk = clk;
    assign pd31_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd31_reset = reset;
    assign pd31_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke_done_out & par0_go_out;
    assign pd32_clk = clk;
    assign pd32_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke0_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd32_reset = reset;
    assign pd32_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke0_done_out & par0_go_out;
    assign pd33_clk = clk;
    assign pd33_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke1_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd33_reset = reset;
    assign pd33_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke1_done_out & par0_go_out;
    assign pd34_clk = clk;
    assign pd34_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke2_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd34_reset = reset;
    assign pd34_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke2_done_out & par0_go_out;
    assign pd35_clk = clk;
    assign pd35_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke3_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd35_reset = reset;
    assign pd35_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke3_done_out & par0_go_out;
    assign pd36_clk = clk;
    assign pd36_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke4_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd36_reset = reset;
    assign pd36_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke4_done_out & par0_go_out;
    assign pd37_clk = clk;
    assign pd37_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke5_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd37_reset = reset;
    assign pd37_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke5_done_out & par0_go_out;
    assign pd38_clk = clk;
    assign pd38_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke6_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd38_reset = reset;
    assign pd38_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke6_done_out & par0_go_out;
    assign pd39_clk = clk;
    assign pd39_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke7_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd39_reset = reset;
    assign pd39_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke7_done_out & par0_go_out;
    assign pd4_clk = clk;
    assign pd4_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc4_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd4_reset = reset;
    assign pd4_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc4_done_out & par_go_out;
    assign pd40_clk = clk;
    assign pd40_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke8_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd40_reset = reset;
    assign pd40_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke8_done_out & par0_go_out;
    assign pd41_clk = clk;
    assign pd41_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke9_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd41_reset = reset;
    assign pd41_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke9_done_out & par0_go_out;
    assign pd42_clk = clk;
    assign pd42_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke10_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd42_reset = reset;
    assign pd42_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke10_done_out & par0_go_out;
    assign pd43_clk = clk;
    assign pd43_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke11_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd43_reset = reset;
    assign pd43_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke11_done_out & par0_go_out;
    assign pd44_clk = clk;
    assign pd44_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke12_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd44_reset = reset;
    assign pd44_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke12_done_out & par0_go_out;
    assign pd45_clk = clk;
    assign pd45_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke13_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd45_reset = reset;
    assign pd45_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke13_done_out & par0_go_out;
    assign pd46_clk = clk;
    assign pd46_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke14_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd46_reset = reset;
    assign pd46_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke14_done_out & par0_go_out;
    assign pd47_clk = clk;
    assign pd47_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke15_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd47_reset = reset;
    assign pd47_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke15_done_out & par0_go_out;
    assign pd48_clk = clk;
    assign pd48_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke16_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd48_reset = reset;
    assign pd48_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke16_done_out & par0_go_out;
    assign pd49_clk = clk;
    assign pd49_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke17_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd49_reset = reset;
    assign pd49_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke17_done_out & par0_go_out;
    assign pd5_clk = clk;
    assign pd5_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc5_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd5_reset = reset;
    assign pd5_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc5_done_out & par_go_out;
    assign pd50_clk = clk;
    assign pd50_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke18_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd50_reset = reset;
    assign pd50_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke18_done_out & par0_go_out;
    assign pd51_clk = clk;
    assign pd51_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke19_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd51_reset = reset;
    assign pd51_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke19_done_out & par0_go_out;
    assign pd52_clk = clk;
    assign pd52_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke20_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd52_reset = reset;
    assign pd52_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke20_done_out & par0_go_out;
    assign pd53_clk = clk;
    assign pd53_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke21_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd53_reset = reset;
    assign pd53_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke21_done_out & par0_go_out;
    assign pd54_clk = clk;
    assign pd54_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke22_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd54_reset = reset;
    assign pd54_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke22_done_out & par0_go_out;
    assign pd55_clk = clk;
    assign pd55_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke23_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd55_reset = reset;
    assign pd55_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke23_done_out & par0_go_out;
    assign pd56_clk = clk;
    assign pd56_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke24_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd56_reset = reset;
    assign pd56_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke24_done_out & par0_go_out;
    assign pd57_clk = clk;
    assign pd57_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke25_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd57_reset = reset;
    assign pd57_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke25_done_out & par0_go_out;
    assign pd58_clk = clk;
    assign pd58_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke26_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd58_reset = reset;
    assign pd58_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke26_done_out & par0_go_out;
    assign pd59_clk = clk;
    assign pd59_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke27_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd59_reset = reset;
    assign pd59_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke27_done_out & par0_go_out;
    assign pd6_clk = clk;
    assign pd6_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc6_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd6_reset = reset;
    assign pd6_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc6_done_out & par_go_out;
    assign pd60_clk = clk;
    assign pd60_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke28_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd60_reset = reset;
    assign pd60_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke28_done_out & par0_go_out;
    assign pd61_clk = clk;
    assign pd61_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke29_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd61_reset = reset;
    assign pd61_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke29_done_out & par0_go_out;
    assign pd62_clk = clk;
    assign pd62_in =
     pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out ? 1'd0 :
     invoke30_done_out & par0_go_out ? 1'd1 : 1'd0;
    assign pd62_reset = reset;
    assign pd62_write_en = pd31_out & pd32_out & pd33_out & pd34_out & pd35_out & pd36_out & pd37_out & pd38_out & pd39_out & pd40_out & pd41_out & pd42_out & pd43_out & pd44_out & pd45_out & pd46_out & pd47_out & pd48_out & pd49_out & pd50_out & pd51_out & pd52_out & pd53_out & pd54_out & pd55_out & pd56_out & pd57_out & pd58_out & pd59_out & pd60_out & pd61_out & pd62_out | invoke30_done_out & par0_go_out;
    assign pd63_clk = clk;
    assign pd63_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke31_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd63_reset = reset;
    assign pd63_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke31_done_out & par1_go_out;
    assign pd64_clk = clk;
    assign pd64_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke32_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd64_reset = reset;
    assign pd64_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke32_done_out & par1_go_out;
    assign pd65_clk = clk;
    assign pd65_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke33_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd65_reset = reset;
    assign pd65_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke33_done_out & par1_go_out;
    assign pd66_clk = clk;
    assign pd66_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke34_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd66_reset = reset;
    assign pd66_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke34_done_out & par1_go_out;
    assign pd67_clk = clk;
    assign pd67_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke35_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd67_reset = reset;
    assign pd67_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke35_done_out & par1_go_out;
    assign pd68_clk = clk;
    assign pd68_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke36_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd68_reset = reset;
    assign pd68_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke36_done_out & par1_go_out;
    assign pd69_clk = clk;
    assign pd69_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke37_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd69_reset = reset;
    assign pd69_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke37_done_out & par1_go_out;
    assign pd7_clk = clk;
    assign pd7_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc7_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd7_reset = reset;
    assign pd7_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc7_done_out & par_go_out;
    assign pd70_clk = clk;
    assign pd70_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke38_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd70_reset = reset;
    assign pd70_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke38_done_out & par1_go_out;
    assign pd71_clk = clk;
    assign pd71_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke39_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd71_reset = reset;
    assign pd71_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke39_done_out & par1_go_out;
    assign pd72_clk = clk;
    assign pd72_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke40_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd72_reset = reset;
    assign pd72_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke40_done_out & par1_go_out;
    assign pd73_clk = clk;
    assign pd73_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke41_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd73_reset = reset;
    assign pd73_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke41_done_out & par1_go_out;
    assign pd74_clk = clk;
    assign pd74_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke42_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd74_reset = reset;
    assign pd74_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke42_done_out & par1_go_out;
    assign pd75_clk = clk;
    assign pd75_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke43_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd75_reset = reset;
    assign pd75_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke43_done_out & par1_go_out;
    assign pd76_clk = clk;
    assign pd76_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke44_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd76_reset = reset;
    assign pd76_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke44_done_out & par1_go_out;
    assign pd77_clk = clk;
    assign pd77_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke45_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd77_reset = reset;
    assign pd77_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke45_done_out & par1_go_out;
    assign pd78_clk = clk;
    assign pd78_in =
     pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out ? 1'd0 :
     invoke46_done_out & par1_go_out ? 1'd1 : 1'd0;
    assign pd78_reset = reset;
    assign pd78_write_en = pd63_out & pd64_out & pd65_out & pd66_out & pd67_out & pd68_out & pd69_out & pd70_out & pd71_out & pd72_out & pd73_out & pd74_out & pd75_out & pd76_out & pd77_out & pd78_out | invoke46_done_out & par1_go_out;
    assign pd79_clk = clk;
    assign pd79_in =
     pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out ? 1'd0 :
     invoke47_done_out & par2_go_out ? 1'd1 : 1'd0;
    assign pd79_reset = reset;
    assign pd79_write_en = pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out | invoke47_done_out & par2_go_out;
    assign pd8_clk = clk;
    assign pd8_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc8_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd8_reset = reset;
    assign pd8_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc8_done_out & par_go_out;
    assign pd80_clk = clk;
    assign pd80_in =
     pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out ? 1'd0 :
     invoke48_done_out & par2_go_out ? 1'd1 : 1'd0;
    assign pd80_reset = reset;
    assign pd80_write_en = pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out | invoke48_done_out & par2_go_out;
    assign pd81_clk = clk;
    assign pd81_in =
     pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out ? 1'd0 :
     invoke49_done_out & par2_go_out ? 1'd1 : 1'd0;
    assign pd81_reset = reset;
    assign pd81_write_en = pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out | invoke49_done_out & par2_go_out;
    assign pd82_clk = clk;
    assign pd82_in =
     pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out ? 1'd0 :
     invoke50_done_out & par2_go_out ? 1'd1 : 1'd0;
    assign pd82_reset = reset;
    assign pd82_write_en = pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out | invoke50_done_out & par2_go_out;
    assign pd83_clk = clk;
    assign pd83_in =
     pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out ? 1'd0 :
     invoke51_done_out & par2_go_out ? 1'd1 : 1'd0;
    assign pd83_reset = reset;
    assign pd83_write_en = pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out | invoke51_done_out & par2_go_out;
    assign pd84_clk = clk;
    assign pd84_in =
     pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out ? 1'd0 :
     invoke52_done_out & par2_go_out ? 1'd1 : 1'd0;
    assign pd84_reset = reset;
    assign pd84_write_en = pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out | invoke52_done_out & par2_go_out;
    assign pd85_clk = clk;
    assign pd85_in =
     pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out ? 1'd0 :
     invoke53_done_out & par2_go_out ? 1'd1 : 1'd0;
    assign pd85_reset = reset;
    assign pd85_write_en = pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out | invoke53_done_out & par2_go_out;
    assign pd86_clk = clk;
    assign pd86_in =
     pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out ? 1'd0 :
     invoke54_done_out & par2_go_out ? 1'd1 : 1'd0;
    assign pd86_reset = reset;
    assign pd86_write_en = pd79_out & pd80_out & pd81_out & pd82_out & pd83_out & pd84_out & pd85_out & pd86_out | invoke54_done_out & par2_go_out;
    assign pd87_clk = clk;
    assign pd87_in =
     pd87_out & pd88_out & pd89_out & pd90_out ? 1'd0 :
     invoke55_done_out & par3_go_out ? 1'd1 : 1'd0;
    assign pd87_reset = reset;
    assign pd87_write_en = pd87_out & pd88_out & pd89_out & pd90_out | invoke55_done_out & par3_go_out;
    assign pd88_clk = clk;
    assign pd88_in =
     pd87_out & pd88_out & pd89_out & pd90_out ? 1'd0 :
     invoke56_done_out & par3_go_out ? 1'd1 : 1'd0;
    assign pd88_reset = reset;
    assign pd88_write_en = pd87_out & pd88_out & pd89_out & pd90_out | invoke56_done_out & par3_go_out;
    assign pd89_clk = clk;
    assign pd89_in =
     pd87_out & pd88_out & pd89_out & pd90_out ? 1'd0 :
     invoke57_done_out & par3_go_out ? 1'd1 : 1'd0;
    assign pd89_reset = reset;
    assign pd89_write_en = pd87_out & pd88_out & pd89_out & pd90_out | invoke57_done_out & par3_go_out;
    assign pd9_clk = clk;
    assign pd9_in =
     pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out ? 1'd0 :
     tdcc9_done_out & par_go_out ? 1'd1 : 1'd0;
    assign pd9_reset = reset;
    assign pd9_write_en = pd_out & pd0_out & pd1_out & pd2_out & pd3_out & pd4_out & pd5_out & pd6_out & pd7_out & pd8_out & pd9_out & pd10_out & pd11_out & pd12_out & pd13_out & pd14_out & pd15_out & pd16_out & pd17_out & pd18_out & pd19_out & pd20_out & pd21_out & pd22_out & pd23_out & pd24_out & pd25_out & pd26_out & pd27_out & pd28_out & pd29_out & pd30_out | tdcc9_done_out & par_go_out;
    assign pd90_clk = clk;
    assign pd90_in =
     pd87_out & pd88_out & pd89_out & pd90_out ? 1'd0 :
     invoke58_done_out & par3_go_out ? 1'd1 : 1'd0;
    assign pd90_reset = reset;
    assign pd90_write_en = pd87_out & pd88_out & pd89_out & pd90_out | invoke58_done_out & par3_go_out;
    assign pd91_clk = clk;
    assign pd91_in =
     pd91_out & pd92_out ? 1'd0 :
     invoke59_done_out & par4_go_out ? 1'd1 : 1'd0;
    assign pd91_reset = reset;
    assign pd91_write_en = pd91_out & pd92_out | invoke59_done_out & par4_go_out;
    assign pd92_clk = clk;
    assign pd92_in =
     pd91_out & pd92_out ? 1'd0 :
     invoke60_done_out & par4_go_out ? 1'd1 : 1'd0;
    assign pd92_reset = reset;
    assign pd92_write_en = pd91_out & pd92_out | invoke60_done_out & par4_go_out;
    assign pd93_clk = clk;
    assign pd93_in =
     pd93_out & pd94_out ? 1'd0 :
     tdcc31_done_out & par5_go_out ? 1'd1 : 1'd0;
    assign pd93_reset = reset;
    assign pd93_write_en = pd93_out & pd94_out | tdcc31_done_out & par5_go_out;
    assign pd94_clk = clk;
    assign pd94_in =
     pd93_out & pd94_out ? 1'd0 :
     tdcc32_done_out & par5_go_out ? 1'd1 : 1'd0;
    assign pd94_reset = reset;
    assign pd94_write_en = pd93_out & pd94_out | tdcc32_done_out & par5_go_out;
    assign save_index_done_in = out_done;
    assign save_index_go_in = ~save_index_done_out & fsm32_out == 4'd7 & tdcc32_go_out;
    assign slice_in =
     write0_go_out | write1_go_out | write2_go_out | write3_go_out | write4_go_out | write5_go_out | write6_go_out | write7_go_out | write8_go_out | write9_go_out | write10_go_out | write11_go_out | write12_go_out | write13_go_out | write14_go_out | write15_go_out | write16_go_out | write17_go_out | write18_go_out | write19_go_out | write20_go_out | write21_go_out | write22_go_out | write23_go_out | write24_go_out | write25_go_out | write26_go_out | write27_go_out | write28_go_out | write29_go_out | write30_go_out | write31_go_out ? sub_out : 6'd0;
    assign sub_left =
     write0_go_out | write1_go_out | write2_go_out | write3_go_out | write4_go_out | write5_go_out | write6_go_out | write7_go_out | write8_go_out | write9_go_out | write10_go_out | write11_go_out | write12_go_out | write13_go_out | write14_go_out | write15_go_out | write16_go_out | write17_go_out | write18_go_out | write19_go_out | write20_go_out | write21_go_out | write22_go_out | write23_go_out | write24_go_out | write25_go_out | write26_go_out | write27_go_out | write28_go_out | write29_go_out | write30_go_out | write31_go_out ? prefix_len : 6'd0;
    assign sub_right =
     write0_go_out | write1_go_out | write2_go_out | write3_go_out | write4_go_out | write5_go_out | write6_go_out | write7_go_out | write8_go_out | write9_go_out | write10_go_out | write11_go_out | write12_go_out | write13_go_out | write14_go_out | write15_go_out | write16_go_out | write17_go_out | write18_go_out | write19_go_out | write20_go_out | write21_go_out | write22_go_out | write23_go_out | write24_go_out | write25_go_out | write26_go_out | write27_go_out | write28_go_out | write29_go_out | write30_go_out | write31_go_out ? 6'd1 : 6'd0;
    assign tdcc0_done_in = fsm0_out == 2'd2;
    assign tdcc0_go_in = ~(pd0_out | tdcc0_done_out) & par_go_out;
    assign tdcc10_done_in = fsm10_out == 2'd2;
    assign tdcc10_go_in = ~(pd10_out | tdcc10_done_out) & par_go_out;
    assign tdcc11_done_in = fsm11_out == 2'd2;
    assign tdcc11_go_in = ~(pd11_out | tdcc11_done_out) & par_go_out;
    assign tdcc12_done_in = fsm12_out == 2'd2;
    assign tdcc12_go_in = ~(pd12_out | tdcc12_done_out) & par_go_out;
    assign tdcc13_done_in = fsm13_out == 2'd2;
    assign tdcc13_go_in = ~(pd13_out | tdcc13_done_out) & par_go_out;
    assign tdcc14_done_in = fsm14_out == 2'd2;
    assign tdcc14_go_in = ~(pd14_out | tdcc14_done_out) & par_go_out;
    assign tdcc15_done_in = fsm15_out == 2'd2;
    assign tdcc15_go_in = ~(pd15_out | tdcc15_done_out) & par_go_out;
    assign tdcc16_done_in = fsm16_out == 2'd2;
    assign tdcc16_go_in = ~(pd16_out | tdcc16_done_out) & par_go_out;
    assign tdcc17_done_in = fsm17_out == 2'd2;
    assign tdcc17_go_in = ~(pd17_out | tdcc17_done_out) & par_go_out;
    assign tdcc18_done_in = fsm18_out == 2'd2;
    assign tdcc18_go_in = ~(pd18_out | tdcc18_done_out) & par_go_out;
    assign tdcc19_done_in = fsm19_out == 2'd2;
    assign tdcc19_go_in = ~(pd19_out | tdcc19_done_out) & par_go_out;
    assign tdcc1_done_in = fsm1_out == 2'd2;
    assign tdcc1_go_in = ~(pd1_out | tdcc1_done_out) & par_go_out;
    assign tdcc20_done_in = fsm20_out == 2'd2;
    assign tdcc20_go_in = ~(pd20_out | tdcc20_done_out) & par_go_out;
    assign tdcc21_done_in = fsm21_out == 2'd2;
    assign tdcc21_go_in = ~(pd21_out | tdcc21_done_out) & par_go_out;
    assign tdcc22_done_in = fsm22_out == 2'd2;
    assign tdcc22_go_in = ~(pd22_out | tdcc22_done_out) & par_go_out;
    assign tdcc23_done_in = fsm23_out == 2'd2;
    assign tdcc23_go_in = ~(pd23_out | tdcc23_done_out) & par_go_out;
    assign tdcc24_done_in = fsm24_out == 2'd2;
    assign tdcc24_go_in = ~(pd24_out | tdcc24_done_out) & par_go_out;
    assign tdcc25_done_in = fsm25_out == 2'd2;
    assign tdcc25_go_in = ~(pd25_out | tdcc25_done_out) & par_go_out;
    assign tdcc26_done_in = fsm26_out == 2'd2;
    assign tdcc26_go_in = ~(pd26_out | tdcc26_done_out) & par_go_out;
    assign tdcc27_done_in = fsm27_out == 2'd2;
    assign tdcc27_go_in = ~(pd27_out | tdcc27_done_out) & par_go_out;
    assign tdcc28_done_in = fsm28_out == 2'd2;
    assign tdcc28_go_in = ~(pd28_out | tdcc28_done_out) & par_go_out;
    assign tdcc29_done_in = fsm29_out == 2'd2;
    assign tdcc29_go_in = ~(pd29_out | tdcc29_done_out) & par_go_out;
    assign tdcc2_done_in = fsm2_out == 2'd2;
    assign tdcc2_go_in = ~(pd2_out | tdcc2_done_out) & par_go_out;
    assign tdcc30_done_in = fsm30_out == 2'd2;
    assign tdcc30_go_in = ~(pd30_out | tdcc30_done_out) & par_go_out;
    assign tdcc31_done_in = fsm31_out == 3'd5;
    assign tdcc31_go_in = ~(pd93_out | tdcc31_done_out) & par5_go_out;
    assign tdcc32_done_in = fsm32_out == 4'd9;
    assign tdcc32_go_in = ~(pd94_out | tdcc32_done_out) & par5_go_out;
    assign tdcc33_done_in = fsm33_out == 1'd1;
    assign tdcc33_go_in = go;
    assign tdcc3_done_in = fsm3_out == 2'd2;
    assign tdcc3_go_in = ~(pd3_out | tdcc3_done_out) & par_go_out;
    assign tdcc4_done_in = fsm4_out == 2'd2;
    assign tdcc4_go_in = ~(pd4_out | tdcc4_done_out) & par_go_out;
    assign tdcc5_done_in = fsm5_out == 2'd2;
    assign tdcc5_go_in = ~(pd5_out | tdcc5_done_out) & par_go_out;
    assign tdcc6_done_in = fsm6_out == 2'd2;
    assign tdcc6_go_in = ~(pd6_out | tdcc6_done_out) & par_go_out;
    assign tdcc7_done_in = fsm7_out == 2'd2;
    assign tdcc7_go_in = ~(pd7_out | tdcc7_done_out) & par_go_out;
    assign tdcc8_done_in = fsm8_out == 2'd2;
    assign tdcc8_go_in = ~(pd8_out | tdcc8_done_out) & par_go_out;
    assign tdcc9_done_in = fsm9_out == 2'd2;
    assign tdcc9_go_in = ~(pd9_out | tdcc9_done_out) & par_go_out;
    assign tdcc_done_in = fsm_out == 2'd2;
    assign tdcc_go_in = ~(pd_out | tdcc_done_out) & par_go_out;
    assign write0_done_in = p0_done & l0_done;
    assign write0_go_in = ~write0_done_out & fsm_out == 2'd1 & tdcc_go_out;
    assign write10_done_in = p10_done & l10_done;
    assign write10_go_in = ~write10_done_out & fsm9_out == 2'd1 & tdcc9_go_out;
    assign write11_done_in = p11_done & l11_done;
    assign write11_go_in = ~write11_done_out & fsm10_out == 2'd1 & tdcc10_go_out;
    assign write12_done_in = p12_done & l12_done;
    assign write12_go_in = ~write12_done_out & fsm11_out == 2'd1 & tdcc11_go_out;
    assign write13_done_in = p13_done & l13_done;
    assign write13_go_in = ~write13_done_out & fsm12_out == 2'd1 & tdcc12_go_out;
    assign write14_done_in = p14_done & l14_done;
    assign write14_go_in = ~write14_done_out & fsm13_out == 2'd1 & tdcc13_go_out;
    assign write15_done_in = p15_done & l15_done;
    assign write15_go_in = ~write15_done_out & fsm14_out == 2'd1 & tdcc14_go_out;
    assign write16_done_in = p16_done & l16_done;
    assign write16_go_in = ~write16_done_out & fsm15_out == 2'd1 & tdcc15_go_out;
    assign write17_done_in = p17_done & l17_done;
    assign write17_go_in = ~write17_done_out & fsm16_out == 2'd1 & tdcc16_go_out;
    assign write18_done_in = p18_done & l18_done;
    assign write18_go_in = ~write18_done_out & fsm17_out == 2'd1 & tdcc17_go_out;
    assign write19_done_in = p19_done & l19_done;
    assign write19_go_in = ~write19_done_out & fsm18_out == 2'd1 & tdcc18_go_out;
    assign write1_done_in = p1_done & l1_done;
    assign write1_go_in = ~write1_done_out & fsm0_out == 2'd1 & tdcc0_go_out;
    assign write20_done_in = p20_done & l20_done;
    assign write20_go_in = ~write20_done_out & fsm19_out == 2'd1 & tdcc19_go_out;
    assign write21_done_in = p21_done & l21_done;
    assign write21_go_in = ~write21_done_out & fsm20_out == 2'd1 & tdcc20_go_out;
    assign write22_done_in = p22_done & l22_done;
    assign write22_go_in = ~write22_done_out & fsm21_out == 2'd1 & tdcc21_go_out;
    assign write23_done_in = p23_done & l23_done;
    assign write23_go_in = ~write23_done_out & fsm22_out == 2'd1 & tdcc22_go_out;
    assign write24_done_in = p24_done & l24_done;
    assign write24_go_in = ~write24_done_out & fsm23_out == 2'd1 & tdcc23_go_out;
    assign write25_done_in = p25_done & l25_done;
    assign write25_go_in = ~write25_done_out & fsm24_out == 2'd1 & tdcc24_go_out;
    assign write26_done_in = p26_done & l26_done;
    assign write26_go_in = ~write26_done_out & fsm25_out == 2'd1 & tdcc25_go_out;
    assign write27_done_in = p27_done & l27_done;
    assign write27_go_in = ~write27_done_out & fsm26_out == 2'd1 & tdcc26_go_out;
    assign write28_done_in = p28_done & l28_done;
    assign write28_go_in = ~write28_done_out & fsm27_out == 2'd1 & tdcc27_go_out;
    assign write29_done_in = p29_done & l29_done;
    assign write29_go_in = ~write29_done_out & fsm28_out == 2'd1 & tdcc28_go_out;
    assign write2_done_in = p2_done & l2_done;
    assign write2_go_in = ~write2_done_out & fsm1_out == 2'd1 & tdcc1_go_out;
    assign write30_done_in = p30_done & l30_done;
    assign write30_go_in = ~write30_done_out & fsm29_out == 2'd1 & tdcc29_go_out;
    assign write31_done_in = p31_done & l31_done;
    assign write31_go_in = ~write31_done_out & fsm30_out == 2'd1 & tdcc30_go_out;
    assign write3_done_in = p3_done & l3_done;
    assign write3_go_in = ~write3_done_out & fsm2_out == 2'd1 & tdcc2_go_out;
    assign write4_done_in = p4_done & l4_done;
    assign write4_go_in = ~write4_done_out & fsm3_out == 2'd1 & tdcc3_go_out;
    assign write5_done_in = p5_done & l5_done;
    assign write5_go_in = ~write5_done_out & fsm4_out == 2'd1 & tdcc4_go_out;
    assign write6_done_in = p6_done & l6_done;
    assign write6_go_in = ~write6_done_out & fsm5_out == 2'd1 & tdcc5_go_out;
    assign write7_done_in = p7_done & l7_done;
    assign write7_go_in = ~write7_done_out & fsm6_out == 2'd1 & tdcc6_go_out;
    assign write8_done_in = p8_done & l8_done;
    assign write8_go_in = ~write8_done_out & fsm7_out == 2'd1 & tdcc7_go_out;
    assign write9_done_in = p9_done & l9_done;
    assign write9_go_in = ~write9_done_out & fsm8_out == 2'd1 & tdcc8_go_out;
    assign write_zero_done_in = zero_index_done;
    assign write_zero_go_in = ~write_zero_done_out & fsm31_out == 3'd2 & tdcc31_go_out;
    assign z_eq_left =
     is_length_zero0_go_out ? 6'd0 : 6'd0;
    assign z_eq_right =
     is_length_zero0_go_out ? prefix_len : 6'd0;
    assign zero_index_clk = clk;
    assign zero_index_in =
     write_zero_go_out ? write_index : 5'd0;
    assign zero_index_reset = reset;
    assign zero_index_write_en = write_zero_go_out;
endmodule

