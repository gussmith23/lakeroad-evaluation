module ugt6_2(input unsigned[5:0] a, input unsigned[5:0] b, output unsigned[5:0] out);
  assign out = a > b;
endmodule
