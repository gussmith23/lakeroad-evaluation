module ugt1_2(input unsigned[0:0] a, input unsigned[0:0] b, output unsigned out);
  assign out = a > b;
endmodule
