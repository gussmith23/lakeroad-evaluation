module sgt4_2(input signed [3:0] a, input signed [3:0] b, output signed out);
  assign out = a > b;
endmodule
