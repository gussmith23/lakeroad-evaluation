module example(input [0:0] a, output[0:0] out);
  assign out = ! a;
endmodule
