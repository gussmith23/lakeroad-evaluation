module ult5_2(input unsigned[4:0] a, input unsigned[4:0] b, output unsigned out);
  assign out = a < b;
endmodule
