module divs6_2(input signed[5:0] a, input signed[5:0] b, output signed[5:0] out);
  assign out = a / b;
endmodule
