module icmp_gt16(input [15:0] a, input [15:0] b, output [0:0] out);
  assign out = a > b;
endmodule
