module extract8_4_2(input [7:0] a, output [3:0] out);
  assign out = a[5:2];
endmodule