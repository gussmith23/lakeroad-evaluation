module add1_2(input [0:0] a, input [0:0] b, output [0:0] out);
  assign out = a + b;
endmodule
