module sadd2_2(input signed[1:0] a, input signed[1:0] b, output signed[1:0] out);
  assign out = a + b;
endmodule
