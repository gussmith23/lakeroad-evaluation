module or4_2(input [3:0] a, input [3:0] b, output [3:0] out);
  assign out = a | b;
endmodule
