module not7_1(input  [6:0] a, output [6:0] out);
  assign out = ~a;
endmodule
