(* use_dsp = "yes" *) module mult_0_stage_unsigned_3_bit(
	input  [2:0] a,
	input  [2:0] b,
	output [2:0] out,
	input clk);

	assign out = a * b;
endmodule
