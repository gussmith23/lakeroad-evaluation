module slt16_2(input signed [15:0] a, input signed [15:0] b, output signed out);
  assign out = a < b;
endmodule
