(* use_dsp = "yes" *) module preaddmul_0_stage_signed_15_bit(
	input signed [14:0] d,
	input signed [14:0] a,
	input signed [14:0] b,
	output [14:0] out,
	input clk);

	assign out = (d + a) * b;
endmodule
