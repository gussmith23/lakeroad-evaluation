module example(input [15:0] a, output [15:0] out);
  assign out = ~ a;
endmodule
