module sgt1_2(input signed [0:0] a, input signed [0:0] b, output signed out);
  assign out = a > b;
endmodule
