module uge1_2(input  [0:0] a, input  [0:0] b, output  out);
  assign out = a >= b;
endmodule
