module sub96_2(input  [95:0] a, input  [95:0] b, output [95:0] out);
  assign out = a - b;
endmodule
