module uge4_2(input unsigned[3:0] a, input unsigned[3:0] b, output unsigned out);
  assign out = a >= b;
endmodule
