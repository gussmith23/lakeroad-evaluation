module sub7_2(input  [6:0] a, input  [6:0] b, output [6:0] out);
  assign out = a - b;
endmodule
