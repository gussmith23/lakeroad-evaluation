module uge2_2(input unsigned[1:0] a, input unsigned[1:0] b, output unsigned out);
  assign out = a >= b;
endmodule
