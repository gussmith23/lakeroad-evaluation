(* use_dsp = "yes" *) module addaddsquare_b_1_stage_unsigned_3_bit(
	input  [2:0] b,
	input  [2:0] c,
	input  [2:0] d,
	output [2:0] out,
	input clk);

	logic  [5:0] stage0;

	always @(posedge clk) begin
	stage0 <= c + ((d + b) * (d + b));

	end

	assign out = stage0;
endmodule
