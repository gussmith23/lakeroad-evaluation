module slt7_2(input signed[6:0] a, input signed[6:0] b, output signed out);
  assign out = a < b;
endmodule
