module icmp_gt8(input [7:0] a, input [7:0] b, output [0:0] out);
  assign out = a > b;
endmodule
