module not64_1(input [63:0] a, output [63:0] out);
  assign out = ~a;
endmodule
