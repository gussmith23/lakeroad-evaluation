module uge6_2(input  [5:0] a, input  [5:0] b, output  out);
  assign out = a >= b;
endmodule
