module uge16_2(input  [15:0] a, input  [15:0] b, output  out);
  assign out = a >= b;
endmodule
