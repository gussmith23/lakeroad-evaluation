module slt8_2(input signed[7:0] a, input signed[7:0] b, output signed out);
  assign out = a < b;
endmodule
