module not5_1(input  [4:0] a, output [4:0] out);
  assign out = ~a;
endmodule
