module not3_1(input  [2:0] a, output [2:0] out);
  assign out = ~a;
endmodule
