module ule7_2(input  [6:0] a, input  [6:0] b, output  out);
  assign out = a <= b;
endmodule
