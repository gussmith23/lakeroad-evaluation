module add5_2(input  [4:0] a, input  [4:0] b, output [4:0] out);
  assign out = a + b;
endmodule
