module extract4_3_1(input [3:0] a, output [2:0] out);
  assign out = a[3:1];
endmodule