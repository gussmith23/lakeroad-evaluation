module not6_1(input  [5:0] a, output [5:0] out);
  assign out = ~a;
endmodule
