module ugt32_2(input unsigned[31:0] a, input unsigned[31:0] b, output unsigned out);
  assign out = a > b;
endmodule
