(* use_dsp = "yes" *) module preaddmul_0_stage_unsigned_13_bit(
	input  [12:0] d,
	input  [12:0] a,
	input  [12:0] b,
	output [12:0] out,
	input clk);

	assign out = (d + a) * b;
endmodule
