module example(input [23:0] a, output [23:0] out);
  assign out = ~ a;
endmodule
