module ule64_2(input  [63:0] a, input  [63:0] b, output  out);
  assign out = a <= b;
endmodule
