module ssub3_2(input signed[2:0] a, input signed[2:0] b, output signed[2:0] out);
  assign out = a - b;
endmodule
