module divu1_2(input unsigned[0:0] a, input unsigned[0:0] b, output unsigned[0:0] out);
  assign out = a / b;
endmodule
